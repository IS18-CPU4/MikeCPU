`default_nettype none

module fsqrt
   ( input wire [31:0] x,
     output wire [31:0] y,
     output wire ovf);

   // split sequence to each subsequence
   wire xs;
   wire [7:0] xe;
   wire [22:0] xm;
   assign {xs, xe, xm} = x;

   // calc s
   wire s;
   assign s = xs;

   wire [7:0] shift_xe;
   assign shift_xe = xe >> 1;

   // calc e
   wire [7:0] e;
   assign e = (xe[0] == 1) ? 8'd189 - shift_xe : 8'd190 - shift_xe; 

   // calc m
   wire [22:0] m;
   wire [45:0] val;
   wire [10:0] key;
   assign key = {xe[0], xm[22:13]};
   // lookup table and get constant and grad
   lookup_table lt(key, val);
   wire [22:0] constant;
   wire [22:0] grad;
   // constant supplements 1 at the MSB
   assign constant = val[45:23];
   assign grad = val[22:0];
   wire [45:0] grad2;
   assign grad2 = xm * grad;
   assign m = constant - grad2;

   wire [31:0] tmp_y;
   fmul u1(x, {s, e, m}, tmp_y, ovf);

   wire [31:0] root2;
   assign root2 = 31'b00111111101101010000010011110011;

   wire [7:0] odd_zero_ye;
   assign odd_zero_ye = shift_xe + 8'd64;

   wire [31:0] even_zero_y;
   wire [7:0] even_zero_tmp_ye;
   assign even_zero_y = 8'd63 + shift_xe;
   wire tmp_ovf;
   fmul u2(root2, {xs, even_zero_tmp_ye, xm}, even_zero_y, tmp_ovf);

   assign y = (xm != 23'd0) ? tmp_y :
              (xe[0] == 1) ? {xs, odd_zero_ye, xm} : even_zero_y;

endmodule

module lookup_table
   ( input wire [10:0] key,
     output wire [45:0] value);

   assign value =
(key == 11'b00000000000) ? 46'b0111111111101000000001001111111111010000000010 :
(key == 11'b00000000001) ? 46'b0111111110111000000101101111111101110000001011 :
(key == 11'b00000000010) ? 46'b0111111110001000001110101111111100010000011101 :
(key == 11'b00000000011) ? 46'b0111111101011000011100001111111010110000111000 :
(key == 11'b00000000100) ? 46'b0111111100101000101110001111111001010001011100 :
(key == 11'b00000000101) ? 46'b0111111011111001000100001111110111110010001000 :
(key == 11'b00000000110) ? 46'b0111111011001001011111001111110110010010111110 :
(key == 11'b00000000111) ? 46'b0111111010011001111111001111110100110011111110 :
(key == 11'b00000001000) ? 46'b0111111001101010100010001111110011010101000100 :
(key == 11'b00000001001) ? 46'b0111111000111011001010101111110001110110010101 :
(key == 11'b00000001010) ? 46'b0111111000001011110111001111110000010111101110 :
(key == 11'b00000001011) ? 46'b0111110111011100100111001111101110111001001110 :
(key == 11'b00000001100) ? 46'b0111110110101101011101001111101101011010111010 :
(key == 11'b00000001101) ? 46'b0111110101111110010110101111101011111100101101 :
(key == 11'b00000001110) ? 46'b0111110101001111010100001111101010011110101000 :
(key == 11'b00000001111) ? 46'b0111110100100000010110001111101001000000101100 :
(key == 11'b00000010000) ? 46'b0111110011110001011101001111100111100010111010 :
(key == 11'b00000010001) ? 46'b0111110011000010101000001111100110000101010000 :
(key == 11'b00000010010) ? 46'b0111110010010011110111101111100100100111101111 :
(key == 11'b00000010011) ? 46'b0111110001100101001011001111100011001010010110 :
(key == 11'b00000010100) ? 46'b0111110000110110100011001111100001101101000110 :
(key == 11'b00000010101) ? 46'b0111110000000111111111001111100000001111111110 :
(key == 11'b00000010110) ? 46'b0111101111011001011111001111011110110010111110 :
(key == 11'b00000010111) ? 46'b0111101110101011000011101111011101010110000111 :
(key == 11'b00000011000) ? 46'b0111101101111100101100101111011011111001011001 :
(key == 11'b00000011001) ? 46'b0111101101001110011010001111011010011100110100 :
(key == 11'b00000011010) ? 46'b0111101100100000001011101111011001000000010111 :
(key == 11'b00000011011) ? 46'b0111101011110010000001001111010111100100000010 :
(key == 11'b00000011100) ? 46'b0111101011000011111010101111010110000111110101 :
(key == 11'b00000011101) ? 46'b0111101010010101111000101111010100101011110001 :
(key == 11'b00000011110) ? 46'b0111101001100111111011001111010011001111110110 :
(key == 11'b00000011111) ? 46'b0111101000111010000001001111010001110100000010 :
(key == 11'b00000100000) ? 46'b0111101000001100001100001111010000011000011000 :
(key == 11'b00000100001) ? 46'b0111100111011110011010101111001110111100110101 :
(key == 11'b00000100010) ? 46'b0111100110110000101101101111001101100001011011 :
(key == 11'b00000100011) ? 46'b0111100110000011000101001111001100000110001010 :
(key == 11'b00000100100) ? 46'b0111100101010101100000001111001010101011000000 :
(key == 11'b00000100101) ? 46'b0111100100100111111111001111001001001111111110 :
(key == 11'b00000100110) ? 46'b0111100011111010100011001111000111110101000110 :
(key == 11'b00000100111) ? 46'b0111100011001101001010001111000110011010010100 :
(key == 11'b00000101000) ? 46'b0111100010011111110101101111000100111111101011 :
(key == 11'b00000101001) ? 46'b0111100001110010100101001111000011100101001010 :
(key == 11'b00000101010) ? 46'b0111100001000101011001001111000010001010110010 :
(key == 11'b00000101011) ? 46'b0111100000011000010000001111000000110000100000 :
(key == 11'b00000101100) ? 46'b0111011111101011001100101110111111010110011001 :
(key == 11'b00000101101) ? 46'b0111011110111110001100101110111101111100011001 :
(key == 11'b00000101110) ? 46'b0111011110010001010000101110111100100010100001 :
(key == 11'b00000101111) ? 46'b0111011101100100011000101110111011001000110001 :
(key == 11'b00000110000) ? 46'b0111011100110111100100101110111001101111001001 :
(key == 11'b00000110001) ? 46'b0111011100001010110100001110111000010101101000 :
(key == 11'b00000110010) ? 46'b0111011011011110001000101110110110111100010001 :
(key == 11'b00000110011) ? 46'b0111011010110001100000101110110101100011000001 :
(key == 11'b00000110100) ? 46'b0111011010000100111100001110110100001001111000 :
(key == 11'b00000110101) ? 46'b0111011001011000011100101110110010110000111001 :
(key == 11'b00000110110) ? 46'b0111011000101100000000101110110001011000000001 :
(key == 11'b00000110111) ? 46'b0111010111111111101000001110101111111111010000 :
(key == 11'b00000111000) ? 46'b0111010111010011010100001110101110100110101000 :
(key == 11'b00000111001) ? 46'b0111010110100111000100001110101101001110001000 :
(key == 11'b00000111010) ? 46'b0111010101111010110111101110101011110101101111 :
(key == 11'b00000111011) ? 46'b0111010101001110101111001110101010011101011110 :
(key == 11'b00000111100) ? 46'b0111010100100010101010001110101001000101010100 :
(key == 11'b00000111101) ? 46'b0111010011110110101010001110100111101101010100 :
(key == 11'b00000111110) ? 46'b0111010011001010101101001110100110010101011010 :
(key == 11'b00000111111) ? 46'b0111010010011110110100101110100100111101101001 :
(key == 11'b00001000000) ? 46'b0111010001110011000000001110100011100110000000 :
(key == 11'b00001000001) ? 46'b0111010001000111001110101110100010001110011101 :
(key == 11'b00001000010) ? 46'b0111010000011011100001001110100000110111000010 :
(key == 11'b00001000011) ? 46'b0111001111101111111000001110011111011111110000 :
(key == 11'b00001000100) ? 46'b0111001111000100010010001110011110001000100100 :
(key == 11'b00001000101) ? 46'b0111001110011000110000001110011100110001100000 :
(key == 11'b00001000110) ? 46'b0111001101101101010010001110011011011010100100 :
(key == 11'b00001000111) ? 46'b0111001101000001111000001110011010000011110000 :
(key == 11'b00001001000) ? 46'b0111001100010110100010001110011000101101000100 :
(key == 11'b00001001001) ? 46'b0111001011101011001111101110010111010110011111 :
(key == 11'b00001001010) ? 46'b0111001011000000000001001110010110000000000010 :
(key == 11'b00001001011) ? 46'b0111001010010100110101101110010100101001101011 :
(key == 11'b00001001100) ? 46'b0111001001101001101110001110010011010011011100 :
(key == 11'b00001001101) ? 46'b0111001000111110101011001110010001111101010110 :
(key == 11'b00001001110) ? 46'b0111001000010011101011101110010000100111010111 :
(key == 11'b00001001111) ? 46'b0111000111101000101111101110001111010001011111 :
(key == 11'b00001010000) ? 46'b0111000110111101110111101110001101111011101111 :
(key == 11'b00001010001) ? 46'b0111000110010011000011001110001100100110000110 :
(key == 11'b00001010010) ? 46'b0111000101101000010010001110001011010000100100 :
(key == 11'b00001010011) ? 46'b0111000100111101100101001110001001111011001010 :
(key == 11'b00001010100) ? 46'b0111000100010010111011101110001000100101110111 :
(key == 11'b00001010101) ? 46'b0111000011101000010110001110000111010000101100 :
(key == 11'b00001010110) ? 46'b0111000010111101110100001110000101111011101000 :
(key == 11'b00001010111) ? 46'b0111000010010011010101101110000100100110101011 :
(key == 11'b00001011000) ? 46'b0111000001101000111011001110000011010001110110 :
(key == 11'b00001011001) ? 46'b0111000000111110100100001110000001111101001000 :
(key == 11'b00001011010) ? 46'b0111000000010100010000001110000000101000100000 :
(key == 11'b00001011011) ? 46'b0110111111101010000001001101111111010100000010 :
(key == 11'b00001011100) ? 46'b0110111110111111110101001101111101111111101010 :
(key == 11'b00001011101) ? 46'b0110111110010101101100001101111100101011011000 :
(key == 11'b00001011110) ? 46'b0110111101101011100111101101111011010111001111 :
(key == 11'b00001011111) ? 46'b0110111101000001100110001101111010000011001100 :
(key == 11'b00001100000) ? 46'b0110111100010111101000101101111000101111010001 :
(key == 11'b00001100001) ? 46'b0110111011101101101110101101110111011011011101 :
(key == 11'b00001100010) ? 46'b0110111011000011111000001101110110000111110000 :
(key == 11'b00001100011) ? 46'b0110111010011010000101101101110100110100001011 :
(key == 11'b00001100100) ? 46'b0110111001110000010110001101110011100000101100 :
(key == 11'b00001100101) ? 46'b0110111001000110101010101101110010001101010101 :
(key == 11'b00001100110) ? 46'b0110111000011101000010001101110000111010000100 :
(key == 11'b00001100111) ? 46'b0110110111110011011101101101101111100110111011 :
(key == 11'b00001101000) ? 46'b0110110111001001111100001101101110010011111000 :
(key == 11'b00001101001) ? 46'b0110110110100000011111001101101101000000111110 :
(key == 11'b00001101010) ? 46'b0110110101110111000101001101101011101110001010 :
(key == 11'b00001101011) ? 46'b0110110101001101101110001101101010011011011100 :
(key == 11'b00001101100) ? 46'b0110110100100100011011001101101001001000110110 :
(key == 11'b00001101101) ? 46'b0110110011111011001100001101100111110110011000 :
(key == 11'b00001101110) ? 46'b0110110011010010000000001101100110100100000000 :
(key == 11'b00001101111) ? 46'b0110110010101000110111001101100101010001101110 :
(key == 11'b00001110000) ? 46'b0110110001111111110010101101100011111111100101 :
(key == 11'b00001110001) ? 46'b0110110001010110110000101101100010101101100001 :
(key == 11'b00001110010) ? 46'b0110110000101101110010001101100001011011100100 :
(key == 11'b00001110011) ? 46'b0110110000000100111000001101100000001001110000 :
(key == 11'b00001110100) ? 46'b0110101111011100000000101101011110111000000001 :
(key == 11'b00001110101) ? 46'b0110101110110011001100001101011101100110011000 :
(key == 11'b00001110110) ? 46'b0110101110001010011100001101011100010100111000 :
(key == 11'b00001110111) ? 46'b0110101101100001101111001101011011000011011110 :
(key == 11'b00001111000) ? 46'b0110101100111001000101001101011001110010001010 :
(key == 11'b00001111001) ? 46'b0110101100010000011111001101011000100000111110 :
(key == 11'b00001111010) ? 46'b0110101011100111111100001101010111001111111000 :
(key == 11'b00001111011) ? 46'b0110101010111111011101001101010101111110111010 :
(key == 11'b00001111100) ? 46'b0110101010010111000001101101010100101110000011 :
(key == 11'b00001111101) ? 46'b0110101001101110101000101101010011011101010001 :
(key == 11'b00001111110) ? 46'b0110101001000110010011101101010010001100100111 :
(key == 11'b00001111111) ? 46'b0110101000011110000010001101010000111100000100 :
(key == 11'b00010000000) ? 46'b0110100111110101110100001101001111101011101000 :
(key == 11'b00010000001) ? 46'b0110100111001101101000001101001110011011010000 :
(key == 11'b00010000010) ? 46'b0110100110100101100000001101001101001011000000 :
(key == 11'b00010000011) ? 46'b0110100101111101011100001101001011111010111000 :
(key == 11'b00010000100) ? 46'b0110100101010101011010101101001010101010110101 :
(key == 11'b00010000101) ? 46'b0110100100101101011101001101001001011010111010 :
(key == 11'b00010000110) ? 46'b0110100100000101100010001101001000001011000100 :
(key == 11'b00010000111) ? 46'b0110100011011101101011001101000110111011010110 :
(key == 11'b00010001000) ? 46'b0110100010110101110111001101000101101011101110 :
(key == 11'b00010001001) ? 46'b0110100010001110000111001101000100011100001110 :
(key == 11'b00010001010) ? 46'b0110100001100110011001001101000011001100110010 :
(key == 11'b00010001011) ? 46'b0110100000111110101111001101000001111101011110 :
(key == 11'b00010001100) ? 46'b0110100000010111001000101101000000101110010001 :
(key == 11'b00010001101) ? 46'b0110011111101111100100101100111111011111001001 :
(key == 11'b00010001110) ? 46'b0110011111001000000100001100111110010000001000 :
(key == 11'b00010001111) ? 46'b0110011110100000101000001100111101000001010000 :
(key == 11'b00010010000) ? 46'b0110011101111001001101101100111011110010011011 :
(key == 11'b00010010001) ? 46'b0110011101010001110111001100111010100011101110 :
(key == 11'b00010010010) ? 46'b0110011100101010100100001100111001010101001000 :
(key == 11'b00010010011) ? 46'b0110011100000011010100001100111000000110101000 :
(key == 11'b00010010100) ? 46'b0110011011011100000111001100110110111000001110 :
(key == 11'b00010010101) ? 46'b0110011010110100111101001100110101101001111010 :
(key == 11'b00010010110) ? 46'b0110011010001101110110101100110100011011101101 :
(key == 11'b00010010111) ? 46'b0110011001100110110011101100110011001101100111 :
(key == 11'b00010011000) ? 46'b0110011000111111110011001100110001111111100110 :
(key == 11'b00010011001) ? 46'b0110011000011000110110001100110000110001101100 :
(key == 11'b00010011010) ? 46'b0110010111110001111100101100101111100011111001 :
(key == 11'b00010011011) ? 46'b0110010111001011000110001100101110010110001100 :
(key == 11'b00010011100) ? 46'b0110010110100100010011001100101101001000100110 :
(key == 11'b00010011101) ? 46'b0110010101111101100011001100101011111011000110 :
(key == 11'b00010011110) ? 46'b0110010101010110110101101100101010101101101011 :
(key == 11'b00010011111) ? 46'b0110010100110000001011001100101001100000010110 :
(key == 11'b00010100000) ? 46'b0110010100001001100101001100101000010011001010 :
(key == 11'b00010100001) ? 46'b0110010011100011000001001100100111000110000010 :
(key == 11'b00010100010) ? 46'b0110010010111100100000101100100101111001000001 :
(key == 11'b00010100011) ? 46'b0110010010010110000011001100100100101100000110 :
(key == 11'b00010100100) ? 46'b0110010001101111101000101100100011011111010001 :
(key == 11'b00010100101) ? 46'b0110010001001001010001001100100010010010100010 :
(key == 11'b00010100110) ? 46'b0110010000100010111101001100100001000101111010 :
(key == 11'b00010100111) ? 46'b0110001111111100101100001100011111111001011000 :
(key == 11'b00010101000) ? 46'b0110001111010110011110001100011110101100111100 :
(key == 11'b00010101001) ? 46'b0110001110110000010011001100011101100000100110 :
(key == 11'b00010101010) ? 46'b0110001110001010001011001100011100010100010110 :
(key == 11'b00010101011) ? 46'b0110001101100100000110001100011011001000001100 :
(key == 11'b00010101100) ? 46'b0110001100111110000100101100011001111100001001 :
(key == 11'b00010101101) ? 46'b0110001100011000000110001100011000110000001100 :
(key == 11'b00010101110) ? 46'b0110001011110010001010001100010111100100010100 :
(key == 11'b00010101111) ? 46'b0110001011001100010001001100010110011000100010 :
(key == 11'b00010110000) ? 46'b0110001010100110011100001100010101001100111000 :
(key == 11'b00010110001) ? 46'b0110001010000000101001101100010100000001010011 :
(key == 11'b00010110010) ? 46'b0110001001011010111010001100010010110101110100 :
(key == 11'b00010110011) ? 46'b0110001000110101001101001100010001101010011010 :
(key == 11'b00010110100) ? 46'b0110001000001111100100001100010000011111001000 :
(key == 11'b00010110101) ? 46'b0110000111101001111101001100001111010011111010 :
(key == 11'b00010110110) ? 46'b0110000111000100011001101100001110001000110011 :
(key == 11'b00010110111) ? 46'b0110000110011110111001101100001100111101110011 :
(key == 11'b00010111000) ? 46'b0110000101111001011100001100001011110010111000 :
(key == 11'b00010111001) ? 46'b0110000101010100000001101100001010101000000011 :
(key == 11'b00010111010) ? 46'b0110000100101110101001001100001001011101010010 :
(key == 11'b00010111011) ? 46'b0110000100001001010100101100001000010010101001 :
(key == 11'b00010111100) ? 46'b0110000011100100000011101100000111001000000111 :
(key == 11'b00010111101) ? 46'b0110000010111110110101001100000101111101101010 :
(key == 11'b00010111110) ? 46'b0110000010011001101000101100000100110011010001 :
(key == 11'b00010111111) ? 46'b0110000001110100011111101100000011101000111111 :
(key == 11'b00011000000) ? 46'b0110000001001111011010001100000010011110110100 :
(key == 11'b00011000001) ? 46'b0110000000101010010110101100000001010100101101 :
(key == 11'b00011000010) ? 46'b0110000000000101010110101100000000001010101101 :
(key == 11'b00011000011) ? 46'b0101111111100000011010001011111111000000110100 :
(key == 11'b00011000100) ? 46'b0101111110111011011111001011111101110110111110 :
(key == 11'b00011000101) ? 46'b0101111110010110101000001011111100101101010000 :
(key == 11'b00011000110) ? 46'b0101111101110001110011001011111011100011100110 :
(key == 11'b00011000111) ? 46'b0101111101001101000010001011111010011010000100 :
(key == 11'b00011001000) ? 46'b0101111100101000010011001011111001010000100110 :
(key == 11'b00011001001) ? 46'b0101111100000011100111001011111000000111001110 :
(key == 11'b00011001010) ? 46'b0101111011011110111110001011110110111101111100 :
(key == 11'b00011001011) ? 46'b0101111010111010011000001011110101110100110000 :
(key == 11'b00011001100) ? 46'b0101111010010101110101001011110100101011101010 :
(key == 11'b00011001101) ? 46'b0101111001110001010100101011110011100010101001 :
(key == 11'b00011001110) ? 46'b0101111001001100110111001011110010011001101110 :
(key == 11'b00011001111) ? 46'b0101111000101000011100101011110001010000111001 :
(key == 11'b00011010000) ? 46'b0101111000000100000100101011110000001000001001 :
(key == 11'b00011010001) ? 46'b0101110111011111101111001011101110111111011110 :
(key == 11'b00011010010) ? 46'b0101110110111011011101001011101101110110111010 :
(key == 11'b00011010011) ? 46'b0101110110010111001110001011101100101110011100 :
(key == 11'b00011010100) ? 46'b0101110101110011000010001011101011100110000100 :
(key == 11'b00011010101) ? 46'b0101110101001110111000001011101010011101110000 :
(key == 11'b00011010110) ? 46'b0101110100101010110000101011101001010101100001 :
(key == 11'b00011010111) ? 46'b0101110100000110101100001011101000001101011000 :
(key == 11'b00011011000) ? 46'b0101110011100010101011001011100111000101010110 :
(key == 11'b00011011001) ? 46'b0101110010111110101101001011100101111101011010 :
(key == 11'b00011011010) ? 46'b0101110010011010110000101011100100110101100001 :
(key == 11'b00011011011) ? 46'b0101110001110110110111001011100011101101101110 :
(key == 11'b00011011100) ? 46'b0101110001010011000001101011100010100110000011 :
(key == 11'b00011011101) ? 46'b0101110000101111001110001011100001011110011100 :
(key == 11'b00011011110) ? 46'b0101110000001011011101101011100000010110111011 :
(key == 11'b00011011111) ? 46'b0101101111100111101111101011011111001111011111 :
(key == 11'b00011100000) ? 46'b0101101111000100000100001011011110001000001000 :
(key == 11'b00011100001) ? 46'b0101101110100000011100001011011101000000111000 :
(key == 11'b00011100010) ? 46'b0101101101111100110101101011011011111001101011 :
(key == 11'b00011100011) ? 46'b0101101101011001010010101011011010110010100101 :
(key == 11'b00011100100) ? 46'b0101101100110101110010101011011001101011100101 :
(key == 11'b00011100101) ? 46'b0101101100010010010101001011011000100100101010 :
(key == 11'b00011100110) ? 46'b0101101011101110111010001011010111011101110100 :
(key == 11'b00011100111) ? 46'b0101101011001011100010001011010110010111000100 :
(key == 11'b00011101000) ? 46'b0101101010101000001100101011010101010000011001 :
(key == 11'b00011101001) ? 46'b0101101010000100111001101011010100001001110011 :
(key == 11'b00011101010) ? 46'b0101101001100001101001101011010011000011010011 :
(key == 11'b00011101011) ? 46'b0101101000111110011100001011010001111100111000 :
(key == 11'b00011101100) ? 46'b0101101000011011010001101011010000110110100011 :
(key == 11'b00011101101) ? 46'b0101100111111000001001001011001111110000010010 :
(key == 11'b00011101110) ? 46'b0101100111010101000100001011001110101010001000 :
(key == 11'b00011101111) ? 46'b0101100110110010000001101011001101100100000011 :
(key == 11'b00011110000) ? 46'b0101100110001111000010001011001100011110000100 :
(key == 11'b00011110001) ? 46'b0101100101101100000100001011001011011000001000 :
(key == 11'b00011110010) ? 46'b0101100101001001001001101011001010010010010011 :
(key == 11'b00011110011) ? 46'b0101100100100110010001101011001001001100100011 :
(key == 11'b00011110100) ? 46'b0101100100000011011100001011001000000110111000 :
(key == 11'b00011110101) ? 46'b0101100011100000101001001011000111000001010010 :
(key == 11'b00011110110) ? 46'b0101100010111101111001001011000101111011110010 :
(key == 11'b00011110111) ? 46'b0101100010011011001011101011000100110110010111 :
(key == 11'b00011111000) ? 46'b0101100001111000100000101011000011110001000001 :
(key == 11'b00011111001) ? 46'b0101100001010101111000001011000010101011110000 :
(key == 11'b00011111010) ? 46'b0101100000110011010010001011000001100110100100 :
(key == 11'b00011111011) ? 46'b0101100000010000101111001011000000100001011110 :
(key == 11'b00011111100) ? 46'b0101011111101110001111001010111111011100011110 :
(key == 11'b00011111101) ? 46'b0101011111001011110001001010111110010111100010 :
(key == 11'b00011111110) ? 46'b0101011110101001010101101010111101010010101011 :
(key == 11'b00011111111) ? 46'b0101011110000110111101001010111100001101111010 :
(key == 11'b00100000000) ? 46'b0101011101100100100110101010111011001001001101 :
(key == 11'b00100000001) ? 46'b0101011101000010010011001010111010000100100110 :
(key == 11'b00100000010) ? 46'b0101011100100000000010001010111001000000000100 :
(key == 11'b00100000011) ? 46'b0101011011111101110100001010110111111011101000 :
(key == 11'b00100000100) ? 46'b0101011011011011101000001010110110110111010000 :
(key == 11'b00100000101) ? 46'b0101011010111001011110001010110101110010111100 :
(key == 11'b00100000110) ? 46'b0101011010010111011000001010110100101110110000 :
(key == 11'b00100000111) ? 46'b0101011001110101010011101010110011101010100111 :
(key == 11'b00100001000) ? 46'b0101011001010011010010001010110010100110100100 :
(key == 11'b00100001001) ? 46'b0101011000110001010011001010110001100010100110 :
(key == 11'b00100001010) ? 46'b0101011000001111010110101010110000011110101101 :
(key == 11'b00100001011) ? 46'b0101010111101101011100001010101111011010111000 :
(key == 11'b00100001100) ? 46'b0101010111001011100100101010101110010111001001 :
(key == 11'b00100001101) ? 46'b0101010110101001101111001010101101010011011110 :
(key == 11'b00100001110) ? 46'b0101010110000111111101001010101100001111111010 :
(key == 11'b00100001111) ? 46'b0101010101100110001101001010101011001100011010 :
(key == 11'b00100010000) ? 46'b0101010101000100011111001010101010001000111110 :
(key == 11'b00100010001) ? 46'b0101010100100010110100001010101001000101101000 :
(key == 11'b00100010010) ? 46'b0101010100000001001011101010101000000010010111 :
(key == 11'b00100010011) ? 46'b0101010011011111100110001010100110111111001100 :
(key == 11'b00100010100) ? 46'b0101010010111110000010001010100101111100000100 :
(key == 11'b00100010101) ? 46'b0101010010011100100001001010100100111001000010 :
(key == 11'b00100010110) ? 46'b0101010001111011000010001010100011110110000100 :
(key == 11'b00100010111) ? 46'b0101010001011001100110001010100010110011001100 :
(key == 11'b00100011000) ? 46'b0101010000111000001100001010100001110000011000 :
(key == 11'b00100011001) ? 46'b0101010000010110110101001010100000101101101010 :
(key == 11'b00100011010) ? 46'b0101001111110101100000001010011111101011000000 :
(key == 11'b00100011011) ? 46'b0101001111010100001110001010011110101000011100 :
(key == 11'b00100011100) ? 46'b0101001110110010111110001010011101100101111100 :
(key == 11'b00100011101) ? 46'b0101001110010001110000001010011100100011100000 :
(key == 11'b00100011110) ? 46'b0101001101110000100101001010011011100001001010 :
(key == 11'b00100011111) ? 46'b0101001101001111011100001010011010011110111000 :
(key == 11'b00100100000) ? 46'b0101001100101110010110001010011001011100101100 :
(key == 11'b00100100001) ? 46'b0101001100001101010010101010011000011010100101 :
(key == 11'b00100100010) ? 46'b0101001011101100010001001010010111011000100010 :
(key == 11'b00100100011) ? 46'b0101001011001011010010001010010110010110100100 :
(key == 11'b00100100100) ? 46'b0101001010101010010101101010010101010100101011 :
(key == 11'b00100100101) ? 46'b0101001010001001011011101010010100010010110111 :
(key == 11'b00100100110) ? 46'b0101001001101000100100001010010011010001001000 :
(key == 11'b00100100111) ? 46'b0101001001000111101110001010010010001111011100 :
(key == 11'b00100101000) ? 46'b0101001000100110111011101010010001001101110111 :
(key == 11'b00100101001) ? 46'b0101001000000110001011001010010000001100010110 :
(key == 11'b00100101010) ? 46'b0101000111100101011101001010001111001010111010 :
(key == 11'b00100101011) ? 46'b0101000111000100110000101010001110001001100001 :
(key == 11'b00100101100) ? 46'b0101000110100100000111001010001101001000001110 :
(key == 11'b00100101101) ? 46'b0101000110000011011111101010001100000110111111 :
(key == 11'b00100101110) ? 46'b0101000101100010111011001010001011000101110110 :
(key == 11'b00100101111) ? 46'b0101000101000010011000101010001010000100110001 :
(key == 11'b00100110000) ? 46'b0101000100100001111001001010001001000011110010 :
(key == 11'b00100110001) ? 46'b0101000100000001011011001010001000000010110110 :
(key == 11'b00100110010) ? 46'b0101000011100000111111101010000111000001111111 :
(key == 11'b00100110011) ? 46'b0101000011000000100111001010000110000001001110 :
(key == 11'b00100110100) ? 46'b0101000010100000010000001010000101000000100000 :
(key == 11'b00100110101) ? 46'b0101000001111111111011101010000011111111110111 :
(key == 11'b00100110110) ? 46'b0101000001011111101001101010000010111111010011 :
(key == 11'b00100110111) ? 46'b0101000000111111011001101010000001111110110011 :
(key == 11'b00100111000) ? 46'b0101000000011111001100101010000000111110011001 :
(key == 11'b00100111001) ? 46'b0100111111111111000001101001111111111110000011 :
(key == 11'b00100111010) ? 46'b0100111111011110111000101001111110111101110001 :
(key == 11'b00100111011) ? 46'b0100111110111110110010001001111101111101100100 :
(key == 11'b00100111100) ? 46'b0100111110011110101110001001111100111101011100 :
(key == 11'b00100111101) ? 46'b0100111101111110101100001001111011111101011000 :
(key == 11'b00100111110) ? 46'b0100111101011110101100001001111010111101011000 :
(key == 11'b00100111111) ? 46'b0100111100111110101111001001111001111101011110 :
(key == 11'b00101000000) ? 46'b0100111100011110110100001001111000111101101000 :
(key == 11'b00101000001) ? 46'b0100111011111110111011001001110111111101110110 :
(key == 11'b00101000010) ? 46'b0100111011011111000101001001110110111110001010 :
(key == 11'b00101000011) ? 46'b0100111010111111010000101001110101111110100001 :
(key == 11'b00101000100) ? 46'b0100111010011111011110101001110100111110111101 :
(key == 11'b00101000101) ? 46'b0100111001111111101111001001110011111111011110 :
(key == 11'b00101000110) ? 46'b0100111001100000000001101001110011000000000011 :
(key == 11'b00101000111) ? 46'b0100111001000000010110101001110010000000101101 :
(key == 11'b00101001000) ? 46'b0100111000100000101101101001110001000001011011 :
(key == 11'b00101001001) ? 46'b0100111000000001000111001001110000000010001110 :
(key == 11'b00101001010) ? 46'b0100110111100001100010101001101111000011000101 :
(key == 11'b00101001011) ? 46'b0100110111000010000000001001101110000100000000 :
(key == 11'b00101001100) ? 46'b0100110110100010100000001001101101000101000000 :
(key == 11'b00101001101) ? 46'b0100110110000011000010101001101100000110000101 :
(key == 11'b00101001110) ? 46'b0100110101100011100111001001101011000111001110 :
(key == 11'b00101001111) ? 46'b0100110101000100001110001001101010001000011100 :
(key == 11'b00101010000) ? 46'b0100110100100100110111001001101001001001101110 :
(key == 11'b00101010001) ? 46'b0100110100000101100010001001101000001011000100 :
(key == 11'b00101010010) ? 46'b0100110011100110001111001001100111001100011110 :
(key == 11'b00101010011) ? 46'b0100110011000110111110101001100110001101111101 :
(key == 11'b00101010100) ? 46'b0100110010100111110000101001100101001111100001 :
(key == 11'b00101010101) ? 46'b0100110010001000100100101001100100010001001001 :
(key == 11'b00101010110) ? 46'b0100110001101001011010101001100011010010110101 :
(key == 11'b00101010111) ? 46'b0100110001001010010011001001100010010100100110 :
(key == 11'b00101011000) ? 46'b0100110000101011001101101001100001010110011011 :
(key == 11'b00101011001) ? 46'b0100110000001100001010001001100000011000010100 :
(key == 11'b00101011010) ? 46'b0100101111101101001001001001011111011010010010 :
(key == 11'b00101011011) ? 46'b0100101111001110001010001001011110011100010100 :
(key == 11'b00101011100) ? 46'b0100101110101111001101001001011101011110011010 :
(key == 11'b00101011101) ? 46'b0100101110010000010010101001011100100000100101 :
(key == 11'b00101011110) ? 46'b0100101101110001011010001001011011100010110100 :
(key == 11'b00101011111) ? 46'b0100101101010010100011101001011010100101000111 :
(key == 11'b00101100000) ? 46'b0100101100110011110000001001011001100111100000 :
(key == 11'b00101100001) ? 46'b0100101100010100111101101001011000101001111011 :
(key == 11'b00101100010) ? 46'b0100101011110110001110001001010111101100011100 :
(key == 11'b00101100011) ? 46'b0100101011010111100000101001010110101111000001 :
(key == 11'b00101100100) ? 46'b0100101010111000110100101001010101110001101001 :
(key == 11'b00101100101) ? 46'b0100101010011010001011001001010100110100010110 :
(key == 11'b00101100110) ? 46'b0100101001111011100011001001010011110111000110 :
(key == 11'b00101100111) ? 46'b0100101001011100111110001001010010111001111100 :
(key == 11'b00101101000) ? 46'b0100101000111110011011001001010001111100110110 :
(key == 11'b00101101001) ? 46'b0100101000011111111010001001010000111111110100 :
(key == 11'b00101101010) ? 46'b0100101000000001011011101001010000000010110111 :
(key == 11'b00101101011) ? 46'b0100100111100010111110101001001111000101111101 :
(key == 11'b00101101100) ? 46'b0100100111000100100100001001001110001001001000 :
(key == 11'b00101101101) ? 46'b0100100110100110001011101001001101001100010111 :
(key == 11'b00101101110) ? 46'b0100100110000111110101001001001100001111101010 :
(key == 11'b00101101111) ? 46'b0100100101101001100000101001001011010011000001 :
(key == 11'b00101110000) ? 46'b0100100101001011001110101001001010010110011101 :
(key == 11'b00101110001) ? 46'b0100100100101100111110101001001001011001111101 :
(key == 11'b00101110010) ? 46'b0100100100001110110000101001001000011101100001 :
(key == 11'b00101110011) ? 46'b0100100011110000100100101001000111100001001001 :
(key == 11'b00101110100) ? 46'b0100100011010010011010001001000110100100110100 :
(key == 11'b00101110101) ? 46'b0100100010110100010010001001000101101000100100 :
(key == 11'b00101110110) ? 46'b0100100010010110001100101001000100101100011001 :
(key == 11'b00101110111) ? 46'b0100100001111000001001001001000011110000010010 :
(key == 11'b00101111000) ? 46'b0100100001011010000111001001000010110100001110 :
(key == 11'b00101111001) ? 46'b0100100000111100000111101001000001111000001111 :
(key == 11'b00101111010) ? 46'b0100100000011110001010001001000000111100010100 :
(key == 11'b00101111011) ? 46'b0100100000000000001110101001000000000000011101 :
(key == 11'b00101111100) ? 46'b0100011111100010010101001000111111000100101010 :
(key == 11'b00101111101) ? 46'b0100011111000100011110001000111110001000111100 :
(key == 11'b00101111110) ? 46'b0100011110100110101000001000111101001101010000 :
(key == 11'b00101111111) ? 46'b0100011110001000110101001000111100010001101010 :
(key == 11'b00110000000) ? 46'b0100011101101011000011101000111011010110000111 :
(key == 11'b00110000001) ? 46'b0100011101001101010100101000111010011010101001 :
(key == 11'b00110000010) ? 46'b0100011100101111100111001000111001011111001110 :
(key == 11'b00110000011) ? 46'b0100011100010001111100001000111000100011111000 :
(key == 11'b00110000100) ? 46'b0100011011110100010011001000110111101000100110 :
(key == 11'b00110000101) ? 46'b0100011011010110101011101000110110101101010111 :
(key == 11'b00110000110) ? 46'b0100011010111001000110001000110101110010001100 :
(key == 11'b00110000111) ? 46'b0100011010011011100011001000110100110111000110 :
(key == 11'b00110001000) ? 46'b0100011001111110000010001000110011111100000100 :
(key == 11'b00110001001) ? 46'b0100011001100000100011001000110011000001000110 :
(key == 11'b00110001010) ? 46'b0100011001000011000101001000110010000110001010 :
(key == 11'b00110001011) ? 46'b0100011000100101101010001000110001001011010100 :
(key == 11'b00110001100) ? 46'b0100011000001000010000101000110000010000100001 :
(key == 11'b00110001101) ? 46'b0100010111101010111001101000101111010101110011 :
(key == 11'b00110001110) ? 46'b0100010111001101100100001000101110011011001000 :
(key == 11'b00110001111) ? 46'b0100010110110000010001001000101101100000100010 :
(key == 11'b00110010000) ? 46'b0100010110010011000000001000101100100110000000 :
(key == 11'b00110010001) ? 46'b0100010101110101110000101000101011101011100001 :
(key == 11'b00110010010) ? 46'b0100010101011000100011001000101010110001000110 :
(key == 11'b00110010011) ? 46'b0100010100111011011000001000101001110110110000 :
(key == 11'b00110010100) ? 46'b0100010100011110001110101000101000111100011101 :
(key == 11'b00110010101) ? 46'b0100010100000001000111001000101000000010001110 :
(key == 11'b00110010110) ? 46'b0100010011100100000001101000100111001000000011 :
(key == 11'b00110010111) ? 46'b0100010011000110111110001000100110001101111100 :
(key == 11'b00110011000) ? 46'b0100010010101001111100001000100101010011111000 :
(key == 11'b00110011001) ? 46'b0100010010001100111100001000100100011001111000 :
(key == 11'b00110011010) ? 46'b0100010001101111111111001000100011011111111110 :
(key == 11'b00110011011) ? 46'b0100010001010011000011001000100010100110000110 :
(key == 11'b00110011100) ? 46'b0100010000110110001001001000100001101100010010 :
(key == 11'b00110011101) ? 46'b0100010000011001010001001000100000110010100010 :
(key == 11'b00110011110) ? 46'b0100001111111100011011001000011111111000110110 :
(key == 11'b00110011111) ? 46'b0100001111011111100111001000011110111111001110 :
(key == 11'b00110100000) ? 46'b0100001111000010110101001000011110000101101010 :
(key == 11'b00110100001) ? 46'b0100001110100110000100101000011101001100001001 :
(key == 11'b00110100010) ? 46'b0100001110001001010110001000011100010010101100 :
(key == 11'b00110100011) ? 46'b0100001101101100101010001000011011011001010100 :
(key == 11'b00110100100) ? 46'b0100001101001111111111101000011010011111111111 :
(key == 11'b00110100101) ? 46'b0100001100110011010111001000011001100110101110 :
(key == 11'b00110100110) ? 46'b0100001100010110110000001000011000101101100000 :
(key == 11'b00110100111) ? 46'b0100001011111010001011101000010111110100010111 :
(key == 11'b00110101000) ? 46'b0100001011011101101000101000010110111011010001 :
(key == 11'b00110101001) ? 46'b0100001011000001001000001000010110000010010000 :
(key == 11'b00110101010) ? 46'b0100001010100100101000001000010101001001010000 :
(key == 11'b00110101011) ? 46'b0100001010001000001011001000010100010000010110 :
(key == 11'b00110101100) ? 46'b0100001001101011110000001000010011010111100000 :
(key == 11'b00110101101) ? 46'b0100001001001111010110001000010010011110101100 :
(key == 11'b00110101110) ? 46'b0100001000110010111110001000010001100101111100 :
(key == 11'b00110101111) ? 46'b0100001000010110101001001000010000101101010010 :
(key == 11'b00110110000) ? 46'b0100000111111010010101001000001111110100101010 :
(key == 11'b00110110001) ? 46'b0100000111011110000011001000001110111100000110 :
(key == 11'b00110110010) ? 46'b0100000111000001110011001000001110000011100110 :
(key == 11'b00110110011) ? 46'b0100000110100101100101001000001101001011001010 :
(key == 11'b00110110100) ? 46'b0100000110001001011000001000001100010010110000 :
(key == 11'b00110110101) ? 46'b0100000101101101001101001000001011011010011010 :
(key == 11'b00110110110) ? 46'b0100000101010001000100101000001010100010001001 :
(key == 11'b00110110111) ? 46'b0100000100110100111101101000001001101001111011 :
(key == 11'b00110111000) ? 46'b0100000100011000111000101000001000110001110001 :
(key == 11'b00110111001) ? 46'b0100000011111100110101101000000111111001101011 :
(key == 11'b00110111010) ? 46'b0100000011100000110100001000000111000001101000 :
(key == 11'b00110111011) ? 46'b0100000011000100110100101000000110001001101001 :
(key == 11'b00110111100) ? 46'b0100000010101000110111001000000101010001101110 :
(key == 11'b00110111101) ? 46'b0100000010001100111011001000000100011001110110 :
(key == 11'b00110111110) ? 46'b0100000001110001000001001000000011100010000010 :
(key == 11'b00110111111) ? 46'b0100000001010101001000101000000010101010010001 :
(key == 11'b00111000000) ? 46'b0100000000111001010010001000000001110010100100 :
(key == 11'b00111000001) ? 46'b0100000000011101011110001000000000111010111100 :
(key == 11'b00111000010) ? 46'b0100000000000001101011001000000000000011010110 :
(key == 11'b00111000011) ? 46'b0011111111100101111010000111111111001011110100 :
(key == 11'b00111000100) ? 46'b0011111111001010001011000111111110010100010110 :
(key == 11'b00111000101) ? 46'b0011111110101110011101000111111101011100111010 :
(key == 11'b00111000110) ? 46'b0011111110010010110001100111111100100101100011 :
(key == 11'b00111000111) ? 46'b0011111101110111001000000111111011101110010000 :
(key == 11'b00111001000) ? 46'b0011111101011011100000000111111010110111000000 :
(key == 11'b00111001001) ? 46'b0011111100111111111001100111111001111111110011 :
(key == 11'b00111001010) ? 46'b0011111100100100010101100111111001001000101011 :
(key == 11'b00111001011) ? 46'b0011111100001000110011000111111000010001100110 :
(key == 11'b00111001100) ? 46'b0011111011101101010010000111110111011010100100 :
(key == 11'b00111001101) ? 46'b0011111011010001110010100111110110100011100101 :
(key == 11'b00111001110) ? 46'b0011111010110110010101000111110101101100101010 :
(key == 11'b00111001111) ? 46'b0011111010011010111010000111110100110101110100 :
(key == 11'b00111010000) ? 46'b0011111001111111100000100111110011111111000001 :
(key == 11'b00111010001) ? 46'b0011111001100100001000100111110011001000010001 :
(key == 11'b00111010010) ? 46'b0011111001001000110010000111110010010001100100 :
(key == 11'b00111010011) ? 46'b0011111000101101011110000111110001011010111100 :
(key == 11'b00111010100) ? 46'b0011111000010010001011000111110000100100010110 :
(key == 11'b00111010101) ? 46'b0011110111110110111010000111101111101101110100 :
(key == 11'b00111010110) ? 46'b0011110111011011101011000111101110110111010110 :
(key == 11'b00111010111) ? 46'b0011110111000000011101100111101110000000111011 :
(key == 11'b00111011000) ? 46'b0011110110100101010001100111101101001010100011 :
(key == 11'b00111011001) ? 46'b0011110110001010001000000111101100010100010000 :
(key == 11'b00111011010) ? 46'b0011110101101110111111100111101011011101111111 :
(key == 11'b00111011011) ? 46'b0011110101010011111001000111101010100111110010 :
(key == 11'b00111011100) ? 46'b0011110100111000110100000111101001110001101000 :
(key == 11'b00111011101) ? 46'b0011110100011101110001000111101000111011100010 :
(key == 11'b00111011110) ? 46'b0011110100000010110000000111101000000101100000 :
(key == 11'b00111011111) ? 46'b0011110011100111110000100111100111001111100001 :
(key == 11'b00111100000) ? 46'b0011110011001100110010100111100110011001100101 :
(key == 11'b00111100001) ? 46'b0011110010110001110110100111100101100011101101 :
(key == 11'b00111100010) ? 46'b0011110010010110111100000111100100101101111000 :
(key == 11'b00111100011) ? 46'b0011110001111100000011000111100011111000000110 :
(key == 11'b00111100100) ? 46'b0011110001100001001100000111100011000010011000 :
(key == 11'b00111100101) ? 46'b0011110001000110010111000111100010001100101110 :
(key == 11'b00111100110) ? 46'b0011110000101011100011100111100001010111000111 :
(key == 11'b00111100111) ? 46'b0011110000010000110010000111100000100001100100 :
(key == 11'b00111101000) ? 46'b0011101111110110000001100111011111101100000011 :
(key == 11'b00111101001) ? 46'b0011101111011011010011100111011110110110100111 :
(key == 11'b00111101010) ? 46'b0011101111000000100110000111011110000001001100 :
(key == 11'b00111101011) ? 46'b0011101110100101111011000111011101001011110110 :
(key == 11'b00111101100) ? 46'b0011101110001011010010000111011100010110100100 :
(key == 11'b00111101101) ? 46'b0011101101110000101010000111011011100001010100 :
(key == 11'b00111101110) ? 46'b0011101101010110000100000111011010101100001000 :
(key == 11'b00111101111) ? 46'b0011101100111011100000000111011001110111000000 :
(key == 11'b00111110000) ? 46'b0011101100100000111101000111011001000001111010 :
(key == 11'b00111110001) ? 46'b0011101100000110011100100111011000001100111001 :
(key == 11'b00111110010) ? 46'b0011101011101011111101000111010111010111111010 :
(key == 11'b00111110011) ? 46'b0011101011010001011111100111010110100010111111 :
(key == 11'b00111110100) ? 46'b0011101010110111000011100111010101101110000111 :
(key == 11'b00111110101) ? 46'b0011101010011100101001000111010100111001010010 :
(key == 11'b00111110110) ? 46'b0011101010000010010000100111010100000100100001 :
(key == 11'b00111110111) ? 46'b0011101001100111111001000111010011001111110010 :
(key == 11'b00111111000) ? 46'b0011101001001101100100000111010010011011001000 :
(key == 11'b00111111001) ? 46'b0011101000110011010000100111010001100110100001 :
(key == 11'b00111111010) ? 46'b0011101000011000111110100111010000110001111101 :
(key == 11'b00111111011) ? 46'b0011100111111110101110000111001111111101011100 :
(key == 11'b00111111100) ? 46'b0011100111100100011111000111001111001000111110 :
(key == 11'b00111111101) ? 46'b0011100111001010010010000111001110010100100100 :
(key == 11'b00111111110) ? 46'b0011100110110000000110100111001101100000001101 :
(key == 11'b00111111111) ? 46'b0011100110010101111101000111001100101011111010 :
(key == 11'b01000000000) ? 46'b0011100101111011110100100111001011110111101001 :
(key == 11'b01000000001) ? 46'b0011100101100001101110000111001011000011011100 :
(key == 11'b01000000010) ? 46'b0011100101000111101001000111001010001111010010 :
(key == 11'b01000000011) ? 46'b0011100100101101100110000111001001011011001100 :
(key == 11'b01000000100) ? 46'b0011100100010011100100000111001000100111001000 :
(key == 11'b01000000101) ? 46'b0011100011111001100100000111000111110011001000 :
(key == 11'b01000000110) ? 46'b0011100011011111100101100111000110111111001011 :
(key == 11'b01000000111) ? 46'b0011100011000101101001000111000110001011010010 :
(key == 11'b01000001000) ? 46'b0011100010101011101110000111000101010111011100 :
(key == 11'b01000001001) ? 46'b0011100010010001110100000111000100100011101000 :
(key == 11'b01000001010) ? 46'b0011100001110111111100000111000011101111111000 :
(key == 11'b01000001011) ? 46'b0011100001011110000110000111000010111100001100 :
(key == 11'b01000001100) ? 46'b0011100001000100010001000111000010001000100010 :
(key == 11'b01000001101) ? 46'b0011100000101010011101100111000001010100111011 :
(key == 11'b01000001110) ? 46'b0011100000010000101100000111000000100001011000 :
(key == 11'b01000001111) ? 46'b0011011111110110111100000110111111101101111000 :
(key == 11'b01000010000) ? 46'b0011011111011101001110000110111110111010011100 :
(key == 11'b01000010001) ? 46'b0011011111000011100001000110111110000111000010 :
(key == 11'b01000010010) ? 46'b0011011110101001110110000110111101010011101100 :
(key == 11'b01000010011) ? 46'b0011011110010000001100000110111100100000011000 :
(key == 11'b01000010100) ? 46'b0011011101110110100100000110111011101101001000 :
(key == 11'b01000010101) ? 46'b0011011101011100111101100110111010111001111011 :
(key == 11'b01000010110) ? 46'b0011011101000011011001000110111010000110110010 :
(key == 11'b01000010111) ? 46'b0011011100101001110110000110111001010011101100 :
(key == 11'b01000011000) ? 46'b0011011100010000010100000110111000100000101000 :
(key == 11'b01000011001) ? 46'b0011011011110110110011100110110111101101100111 :
(key == 11'b01000011010) ? 46'b0011011011011101010101000110110110111010101010 :
(key == 11'b01000011011) ? 46'b0011011011000011111000000110110110000111110000 :
(key == 11'b01000011100) ? 46'b0011011010101010011100100110110101010100111001 :
(key == 11'b01000011101) ? 46'b0011011010010001000010000110110100100010000100 :
(key == 11'b01000011110) ? 46'b0011011001110111101010000110110011101111010100 :
(key == 11'b01000011111) ? 46'b0011011001011110010011100110110010111100100111 :
(key == 11'b01000100000) ? 46'b0011011001000100111110000110110010001001111100 :
(key == 11'b01000100001) ? 46'b0011011000101011101010000110110001010111010100 :
(key == 11'b01000100010) ? 46'b0011011000010010011000000110110000100100110000 :
(key == 11'b01000100011) ? 46'b0011010111111001000111100110101111110010001111 :
(key == 11'b01000100100) ? 46'b0011010111011111111000100110101110111111110001 :
(key == 11'b01000100101) ? 46'b0011010111000110101011000110101110001101010110 :
(key == 11'b01000100110) ? 46'b0011010110101101011111000110101101011010111110 :
(key == 11'b01000100111) ? 46'b0011010110010100010100100110101100101000101001 :
(key == 11'b01000101000) ? 46'b0011010101111011001011000110101011110110010110 :
(key == 11'b01000101001) ? 46'b0011010101100010000100000110101011000100001000 :
(key == 11'b01000101010) ? 46'b0011010101001000111110000110101010010001111100 :
(key == 11'b01000101011) ? 46'b0011010100101111111010000110101001011111110100 :
(key == 11'b01000101100) ? 46'b0011010100010110110111000110101000101101101110 :
(key == 11'b01000101101) ? 46'b0011010011111101110101100110100111111011101011 :
(key == 11'b01000101110) ? 46'b0011010011100100110110000110100111001001101100 :
(key == 11'b01000101111) ? 46'b0011010011001011111000000110100110010111110000 :
(key == 11'b01000110000) ? 46'b0011010010110010111011000110100101100101110110 :
(key == 11'b01000110001) ? 46'b0011010010011010000000000110100100110100000000 :
(key == 11'b01000110010) ? 46'b0011010010000001000110000110100100000010001100 :
(key == 11'b01000110011) ? 46'b0011010001101000001110000110100011010000011100 :
(key == 11'b01000110100) ? 46'b0011010001001111010111000110100010011110101110 :
(key == 11'b01000110101) ? 46'b0011010000110110100001100110100001101101000011 :
(key == 11'b01000110110) ? 46'b0011010000011101101110000110100000111011011100 :
(key == 11'b01000110111) ? 46'b0011010000000100111100000110100000001001111000 :
(key == 11'b01000111000) ? 46'b0011001111101100001011000110011111011000010110 :
(key == 11'b01000111001) ? 46'b0011001111010011011100000110011110100110111000 :
(key == 11'b01000111010) ? 46'b0011001110111010101110000110011101110101011100 :
(key == 11'b01000111011) ? 46'b0011001110100010000010000110011101000100000100 :
(key == 11'b01000111100) ? 46'b0011001110001001010111000110011100010010101110 :
(key == 11'b01000111101) ? 46'b0011001101110000101110000110011011100001011100 :
(key == 11'b01000111110) ? 46'b0011001101011000000110000110011010110000001100 :
(key == 11'b01000111111) ? 46'b0011001100111111011111100110011001111110111111 :
(key == 11'b01001000000) ? 46'b0011001100100110111011000110011001001101110110 :
(key == 11'b01001000001) ? 46'b0011001100001110010111000110011000011100101110 :
(key == 11'b01001000010) ? 46'b0011001011110101110101000110010111101011101010 :
(key == 11'b01001000011) ? 46'b0011001011011101010101000110010110111010101010 :
(key == 11'b01001000100) ? 46'b0011001011000100110110000110010110001001101100 :
(key == 11'b01001000101) ? 46'b0011001010101100011000100110010101011000110001 :
(key == 11'b01001000110) ? 46'b0011001010010011111100100110010100100111111001 :
(key == 11'b01001000111) ? 46'b0011001001111011100010000110010011110111000100 :
(key == 11'b01001001000) ? 46'b0011001001100011001000000110010011000110010000 :
(key == 11'b01001001001) ? 46'b0011001001001010110001000110010010010101100010 :
(key == 11'b01001001010) ? 46'b0011001000110010011010100110010001100100110101 :
(key == 11'b01001001011) ? 46'b0011001000011010000110000110010000110100001100 :
(key == 11'b01001001100) ? 46'b0011001000000001110011000110010000000011100110 :
(key == 11'b01001001101) ? 46'b0011000111101001100001000110001111010011000010 :
(key == 11'b01001001110) ? 46'b0011000111010001010000000110001110100010100000 :
(key == 11'b01001001111) ? 46'b0011000110111001000001100110001101110010000011 :
(key == 11'b01001010000) ? 46'b0011000110100000110100000110001101000001101000 :
(key == 11'b01001010001) ? 46'b0011000110001000101000000110001100010001010000 :
(key == 11'b01001010010) ? 46'b0011000101110000011101000110001011100000111010 :
(key == 11'b01001010011) ? 46'b0011000101011000010100000110001010110000101000 :
(key == 11'b01001010100) ? 46'b0011000101000000001100000110001010000000011000 :
(key == 11'b01001010101) ? 46'b0011000100101000000110000110001001010000001100 :
(key == 11'b01001010110) ? 46'b0011000100010000000001000110001000100000000010 :
(key == 11'b01001010111) ? 46'b0011000011110111111101000110000111101111111010 :
(key == 11'b01001011000) ? 46'b0011000011011111111011000110000110111111110110 :
(key == 11'b01001011001) ? 46'b0011000011000111111010100110000110001111110101 :
(key == 11'b01001011010) ? 46'b0011000010101111111011000110000101011111110110 :
(key == 11'b01001011011) ? 46'b0011000010010111111101000110000100101111111010 :
(key == 11'b01001011100) ? 46'b0011000010000000000001000110000100000000000010 :
(key == 11'b01001011101) ? 46'b0011000001101000000101100110000011010000001011 :
(key == 11'b01001011110) ? 46'b0011000001010000001100000110000010100000011000 :
(key == 11'b01001011111) ? 46'b0011000000111000010011100110000001110000100111 :
(key == 11'b01001100000) ? 46'b0011000000100000011100100110000001000000111001 :
(key == 11'b01001100001) ? 46'b0011000000001000100111000110000000010001001110 :
(key == 11'b01001100010) ? 46'b0010111111110000110011000101111111100001100110 :
(key == 11'b01001100011) ? 46'b0010111111011001000000100101111110110010000001 :
(key == 11'b01001100100) ? 46'b0010111111000001001111100101111110000010011111 :
(key == 11'b01001100101) ? 46'b0010111110101001011111000101111101010010111110 :
(key == 11'b01001100110) ? 46'b0010111110010001110001000101111100100011100010 :
(key == 11'b01001100111) ? 46'b0010111101111010000100000101111011110100001000 :
(key == 11'b01001101000) ? 46'b0010111101100010011000000101111011000100110000 :
(key == 11'b01001101001) ? 46'b0010111101001010101110000101111010010101011100 :
(key == 11'b01001101010) ? 46'b0010111100110011000101000101111001100110001010 :
(key == 11'b01001101011) ? 46'b0010111100011011011110000101111000110110111100 :
(key == 11'b01001101100) ? 46'b0010111100000011110111100101111000000111101111 :
(key == 11'b01001101101) ? 46'b0010111011101100010010100101110111011000100101 :
(key == 11'b01001101110) ? 46'b0010111011010100101111000101110110101001011110 :
(key == 11'b01001101111) ? 46'b0010111010111101001101100101110101111010011011 :
(key == 11'b01001110000) ? 46'b0010111010100101101101000101110101001011011010 :
(key == 11'b01001110001) ? 46'b0010111010001110001101100101110100011100011011 :
(key == 11'b01001110010) ? 46'b0010111001110110101111000101110011101101011110 :
(key == 11'b01001110011) ? 46'b0010111001011111010011000101110010111110100110 :
(key == 11'b01001110100) ? 46'b0010111001000111111000000101110010001111110000 :
(key == 11'b01001110101) ? 46'b0010111000110000011110000101110001100000111100 :
(key == 11'b01001110110) ? 46'b0010111000011001000101000101110000110010001010 :
(key == 11'b01001110111) ? 46'b0010111000000001101110000101110000000011011100 :
(key == 11'b01001111000) ? 46'b0010110111101010011000100101101111010100110001 :
(key == 11'b01001111001) ? 46'b0010110111010011000100000101101110100110001000 :
(key == 11'b01001111010) ? 46'b0010110110111011110001000101101101110111100010 :
(key == 11'b01001111011) ? 46'b0010110110100100011111100101101101001000111111 :
(key == 11'b01001111100) ? 46'b0010110110001101001111000101101100011010011110 :
(key == 11'b01001111101) ? 46'b0010110101110110000000000101101011101100000000 :
(key == 11'b01001111110) ? 46'b0010110101011110110010100101101010111101100101 :
(key == 11'b01001111111) ? 46'b0010110101000111100110000101101010001111001100 :
(key == 11'b01010000000) ? 46'b0010110100110000011011000101101001100000110110 :
(key == 11'b01010000001) ? 46'b0010110100011001010001100101101000110010100011 :
(key == 11'b01010000010) ? 46'b0010110100000010001001000101101000000100010010 :
(key == 11'b01010000011) ? 46'b0010110011101011000010000101100111010110000100 :
(key == 11'b01010000100) ? 46'b0010110011010011111100100101100110100111111001 :
(key == 11'b01010000101) ? 46'b0010110010111100111000000101100101111001110000 :
(key == 11'b01010000110) ? 46'b0010110010100101110101000101100101001011101010 :
(key == 11'b01010000111) ? 46'b0010110010001110110011100101100100011101100111 :
(key == 11'b01010001000) ? 46'b0010110001110111110011000101100011101111100110 :
(key == 11'b01010001001) ? 46'b0010110001100000110100000101100011000001101000 :
(key == 11'b01010001010) ? 46'b0010110001001001110110000101100010010011101100 :
(key == 11'b01010001011) ? 46'b0010110000110010111001100101100001100101110011 :
(key == 11'b01010001100) ? 46'b0010110000011011111110100101100000110111111101 :
(key == 11'b01010001101) ? 46'b0010110000000101000101000101100000001010001010 :
(key == 11'b01010001110) ? 46'b0010101111101110001101000101011111011100011010 :
(key == 11'b01010001111) ? 46'b0010101111010111010101100101011110101110101011 :
(key == 11'b01010010000) ? 46'b0010101111000000011111000101011110000000111110 :
(key == 11'b01010010001) ? 46'b0010101110101001101011000101011101010011010110 :
(key == 11'b01010010010) ? 46'b0010101110010010110111100101011100100101101111 :
(key == 11'b01010010011) ? 46'b0010101101111100000101100101011011111000001011 :
(key == 11'b01010010100) ? 46'b0010101101100101010101000101011011001010101010 :
(key == 11'b01010010101) ? 46'b0010101101001110100101100101011010011101001011 :
(key == 11'b01010010110) ? 46'b0010101100110111110111100101011001101111101111 :
(key == 11'b01010010111) ? 46'b0010101100100001001011000101011001000010010110 :
(key == 11'b01010011000) ? 46'b0010101100001010011111000101011000010100111110 :
(key == 11'b01010011001) ? 46'b0010101011110011110101000101010111100111101010 :
(key == 11'b01010011010) ? 46'b0010101011011101001100100101010110111010011001 :
(key == 11'b01010011011) ? 46'b0010101011000110100100100101010110001101001001 :
(key == 11'b01010011100) ? 46'b0010101010101111111110100101010101011111111101 :
(key == 11'b01010011101) ? 46'b0010101010011001011001000101010100110010110010 :
(key == 11'b01010011110) ? 46'b0010101010000010110101100101010100000101101011 :
(key == 11'b01010011111) ? 46'b0010101001101100010011000101010011011000100110 :
(key == 11'b01010100000) ? 46'b0010101001010101110001100101010010101011100011 :
(key == 11'b01010100001) ? 46'b0010101000111111010010000101010001111110100100 :
(key == 11'b01010100010) ? 46'b0010101000101000110011000101010001010001100110 :
(key == 11'b01010100011) ? 46'b0010101000010010010101100101010000100100101011 :
(key == 11'b01010100100) ? 46'b0010100111111011111001000101001111110111110010 :
(key == 11'b01010100101) ? 46'b0010100111100101011110100101001111001010111101 :
(key == 11'b01010100110) ? 46'b0010100111001111000101000101001110011110001010 :
(key == 11'b01010100111) ? 46'b0010100110111000101101000101001101110001011010 :
(key == 11'b01010101000) ? 46'b0010100110100010010110000101001101000100101100 :
(key == 11'b01010101001) ? 46'b0010100110001011111111100101001100010111111111 :
(key == 11'b01010101010) ? 46'b0010100101110101101011000101001011101011010110 :
(key == 11'b01010101011) ? 46'b0010100101011111010111100101001010111110101111 :
(key == 11'b01010101100) ? 46'b0010100101001001000110000101001010010010001100 :
(key == 11'b01010101101) ? 46'b0010100100110010110101000101001001100101101010 :
(key == 11'b01010101110) ? 46'b0010100100011100100101000101001000111001001010 :
(key == 11'b01010101111) ? 46'b0010100100000110010111000101001000001100101110 :
(key == 11'b01010110000) ? 46'b0010100011110000001010000101000111100000010100 :
(key == 11'b01010110001) ? 46'b0010100011011001111110000101000110110011111100 :
(key == 11'b01010110010) ? 46'b0010100011000011110011000101000110000111100110 :
(key == 11'b01010110011) ? 46'b0010100010101101101010000101000101011011010100 :
(key == 11'b01010110100) ? 46'b0010100010010111100010000101000100101111000100 :
(key == 11'b01010110101) ? 46'b0010100010000001011011000101000100000010110110 :
(key == 11'b01010110110) ? 46'b0010100001101011010101100101000011010110101011 :
(key == 11'b01010110111) ? 46'b0010100001010101010001000101000010101010100010 :
(key == 11'b01010111000) ? 46'b0010100000111111001110000101000001111110011100 :
(key == 11'b01010111001) ? 46'b0010100000101001001100000101000001010010011000 :
(key == 11'b01010111010) ? 46'b0010100000010011001011000101000000100110010110 :
(key == 11'b01010111011) ? 46'b0010011111111101001011100100111111111010010111 :
(key == 11'b01010111100) ? 46'b0010011111100111001101100100111111001110011011 :
(key == 11'b01010111101) ? 46'b0010011111010001010000100100111110100010100001 :
(key == 11'b01010111110) ? 46'b0010011110111011010100100100111101110110101001 :
(key == 11'b01010111111) ? 46'b0010011110100101011010000100111101001010110100 :
(key == 11'b01011000000) ? 46'b0010011110001111100001000100111100011111000010 :
(key == 11'b01011000001) ? 46'b0010011101111001101001000100111011110011010010 :
(key == 11'b01011000010) ? 46'b0010011101100011110001000100111011000111100010 :
(key == 11'b01011000011) ? 46'b0010011101001101111011100100111010011011110111 :
(key == 11'b01011000100) ? 46'b0010011100111000000111000100111001110000001110 :
(key == 11'b01011000101) ? 46'b0010011100100010010100000100111001000100101000 :
(key == 11'b01011000110) ? 46'b0010011100001100100010000100111000011001000100 :
(key == 11'b01011000111) ? 46'b0010011011110110110001000100110111101101100010 :
(key == 11'b01011001000) ? 46'b0010011011100001000001000100110111000010000010 :
(key == 11'b01011001001) ? 46'b0010011011001011010010100100110110010110100101 :
(key == 11'b01011001010) ? 46'b0010011010110101100101000100110101101011001010 :
(key == 11'b01011001011) ? 46'b0010011010011111111001000100110100111111110010 :
(key == 11'b01011001100) ? 46'b0010011010001010001110000100110100010100011100 :
(key == 11'b01011001101) ? 46'b0010011001110100100100100100110011101001001001 :
(key == 11'b01011001110) ? 46'b0010011001011110111100000100110010111101111000 :
(key == 11'b01011001111) ? 46'b0010011001001001010101000100110010010010101010 :
(key == 11'b01011010000) ? 46'b0010011000110011101111000100110001100111011110 :
(key == 11'b01011010001) ? 46'b0010011000011110001010000100110000111100010100 :
(key == 11'b01011010010) ? 46'b0010011000001000100110000100110000010001001100 :
(key == 11'b01011010011) ? 46'b0010010111110011000011000100101111100110000110 :
(key == 11'b01011010100) ? 46'b0010010111011101100010000100101110111011000100 :
(key == 11'b01011010101) ? 46'b0010010111001000000010000100101110010000000100 :
(key == 11'b01011010110) ? 46'b0010010110110010100011000100101101100101000110 :
(key == 11'b01011010111) ? 46'b0010010110011101000101000100101100111010001010 :
(key == 11'b01011011000) ? 46'b0010010110000111101000000100101100001111010000 :
(key == 11'b01011011001) ? 46'b0010010101110010001101000100101011100100011010 :
(key == 11'b01011011010) ? 46'b0010010101011100110011000100101010111001100110 :
(key == 11'b01011011011) ? 46'b0010010101000111011001000100101010001110110010 :
(key == 11'b01011011100) ? 46'b0010010100110010000001000100101001100100000010 :
(key == 11'b01011011101) ? 46'b0010010100011100101011000100101000111001010110 :
(key == 11'b01011011110) ? 46'b0010010100000111010101000100101000001110101010 :
(key == 11'b01011011111) ? 46'b0010010011110010000000000100100111100100000000 :
(key == 11'b01011100000) ? 46'b0010010011011100101101000100100110111001011010 :
(key == 11'b01011100001) ? 46'b0010010011000111011010100100100110001110110101 :
(key == 11'b01011100010) ? 46'b0010010010110010001001100100100101100100010011 :
(key == 11'b01011100011) ? 46'b0010010010011100111010000100100100111001110100 :
(key == 11'b01011100100) ? 46'b0010010010000111101011000100100100001111010110 :
(key == 11'b01011100101) ? 46'b0010010001110010011110000100100011100100111100 :
(key == 11'b01011100110) ? 46'b0010010001011101010001000100100010111010100010 :
(key == 11'b01011100111) ? 46'b0010010001001000000110000100100010010000001100 :
(key == 11'b01011101000) ? 46'b0010010000110010111100000100100001100101111000 :
(key == 11'b01011101001) ? 46'b0010010000011101110011000100100000111011100110 :
(key == 11'b01011101010) ? 46'b0010010000001000101011000100100000010001010110 :
(key == 11'b01011101011) ? 46'b0010001111110011100100100100011111100111001001 :
(key == 11'b01011101100) ? 46'b0010001111011110011111000100011110111100111110 :
(key == 11'b01011101101) ? 46'b0010001111001001011010100100011110010010110101 :
(key == 11'b01011101110) ? 46'b0010001110110100010111000100011101101000101110 :
(key == 11'b01011101111) ? 46'b0010001110011111010101100100011100111110101011 :
(key == 11'b01011110000) ? 46'b0010001110001010010100000100011100010100101000 :
(key == 11'b01011110001) ? 46'b0010001101110101010100100100011011101010101001 :
(key == 11'b01011110010) ? 46'b0010001101100000010110000100011011000000101100 :
(key == 11'b01011110011) ? 46'b0010001101001011011001000100011010010110110010 :
(key == 11'b01011110100) ? 46'b0010001100110110011100000100011001101100111000 :
(key == 11'b01011110101) ? 46'b0010001100100001100000100100011001000011000001 :
(key == 11'b01011110110) ? 46'b0010001100001100100110000100011000011001001100 :
(key == 11'b01011110111) ? 46'b0010001011110111101110000100010111101111011100 :
(key == 11'b01011111000) ? 46'b0010001011100010110101100100010111000101101011 :
(key == 11'b01011111001) ? 46'b0010001011001101111110100100010110011011111101 :
(key == 11'b01011111010) ? 46'b0010001010111001001001000100010101110010010010 :
(key == 11'b01011111011) ? 46'b0010001010100100010101000100010101001000101010 :
(key == 11'b01011111100) ? 46'b0010001010001111100001000100010100011111000010 :
(key == 11'b01011111101) ? 46'b0010001001111010101110100100010011110101011101 :
(key == 11'b01011111110) ? 46'b0010001001100101111101000100010011001011111010 :
(key == 11'b01011111111) ? 46'b0010001001010001001110000100010010100010011100 :
(key == 11'b01100000000) ? 46'b0010001000111100011110100100010001111000111101 :
(key == 11'b01100000001) ? 46'b0010001000100111110000100100010001001111100001 :
(key == 11'b01100000010) ? 46'b0010001000010011000100000100010000100110001000 :
(key == 11'b01100000011) ? 46'b0010000111111110011000000100001111111100110000 :
(key == 11'b01100000100) ? 46'b0010000111101001101110000100001111010011011100 :
(key == 11'b01100000101) ? 46'b0010000111010101000100000100001110101010001000 :
(key == 11'b01100000110) ? 46'b0010000111000000011100000100001110000000111000 :
(key == 11'b01100000111) ? 46'b0010000110101011110100100100001101010111101001 :
(key == 11'b01100001000) ? 46'b0010000110010111001110100100001100101110011101 :
(key == 11'b01100001001) ? 46'b0010000110000010101001100100001100000101010011 :
(key == 11'b01100001010) ? 46'b0010000101101110000101100100001011011100001011 :
(key == 11'b01100001011) ? 46'b0010000101011001100010100100001010110011000101 :
(key == 11'b01100001100) ? 46'b0010000101000101000001000100001010001010000010 :
(key == 11'b01100001101) ? 46'b0010000100110000100000000100001001100001000000 :
(key == 11'b01100001110) ? 46'b0010000100011100000000100100001000111000000001 :
(key == 11'b01100001111) ? 46'b0010000100000111100010000100001000001111000100 :
(key == 11'b01100010000) ? 46'b0010000011110011000100100100000111100110001001 :
(key == 11'b01100010001) ? 46'b0010000011011110101000100100000110111101010001 :
(key == 11'b01100010010) ? 46'b0010000011001010001101000100000110010100011010 :
(key == 11'b01100010011) ? 46'b0010000010110101110011000100000101101011100110 :
(key == 11'b01100010100) ? 46'b0010000010100001011010000100000101000010110100 :
(key == 11'b01100010101) ? 46'b0010000010001101000010000100000100011010000100 :
(key == 11'b01100010110) ? 46'b0010000001111000101011000100000011110001010110 :
(key == 11'b01100010111) ? 46'b0010000001100100010101000100000011001000101010 :
(key == 11'b01100011000) ? 46'b0010000001010000000000000100000010100000000000 :
(key == 11'b01100011001) ? 46'b0010000000111011101100100100000001110111011001 :
(key == 11'b01100011010) ? 46'b0010000000100111011010000100000001001110110100 :
(key == 11'b01100011011) ? 46'b0010000000010011001001000100000000100110010010 :
(key == 11'b01100011100) ? 46'b0001111111111110111000100011111111111101110001 :
(key == 11'b01100011101) ? 46'b0001111111101010101001000011111111010101010010 :
(key == 11'b01100011110) ? 46'b0001111111010110011010000011111110101100110100 :
(key == 11'b01100011111) ? 46'b0001111111000010001101000011111110000100011010 :
(key == 11'b01100100000) ? 46'b0001111110101110000001000011111101011100000010 :
(key == 11'b01100100001) ? 46'b0001111110011001110101100011111100110011101011 :
(key == 11'b01100100010) ? 46'b0001111110000101101011100011111100001011010111 :
(key == 11'b01100100011) ? 46'b0001111101110001100010100011111011100011000101 :
(key == 11'b01100100100) ? 46'b0001111101011101011010100011111010111010110101 :
(key == 11'b01100100101) ? 46'b0001111101001001010011100011111010010010100111 :
(key == 11'b01100100110) ? 46'b0001111100110101001110000011111001101010011100 :
(key == 11'b01100100111) ? 46'b0001111100100001001001000011111001000010010010 :
(key == 11'b01100101000) ? 46'b0001111100001101000101000011111000011010001010 :
(key == 11'b01100101001) ? 46'b0001111011111001000011000011110111110010000110 :
(key == 11'b01100101010) ? 46'b0001111011100101000001000011110111001010000010 :
(key == 11'b01100101011) ? 46'b0001111011010001000000100011110110100010000001 :
(key == 11'b01100101100) ? 46'b0001111010111101000001000011110101111010000010 :
(key == 11'b01100101101) ? 46'b0001111010101001000010100011110101010010000101 :
(key == 11'b01100101110) ? 46'b0001111010010101000100100011110100101010001001 :
(key == 11'b01100101111) ? 46'b0001111010000001001000100011110100000010010001 :
(key == 11'b01100110000) ? 46'b0001111001101101001101000011110011011010011010 :
(key == 11'b01100110001) ? 46'b0001111001011001010011000011110010110010100110 :
(key == 11'b01100110010) ? 46'b0001111001000101011001000011110010001010110010 :
(key == 11'b01100110011) ? 46'b0001111000110001100001000011110001100011000010 :
(key == 11'b01100110100) ? 46'b0001111000011101101001100011110000111011010011 :
(key == 11'b01100110101) ? 46'b0001111000001001110011100011110000010011100111 :
(key == 11'b01100110110) ? 46'b0001110111110101111110100011101111101011111101 :
(key == 11'b01100110111) ? 46'b0001110111100010001010000011101111000100010100 :
(key == 11'b01100111000) ? 46'b0001110111001110010111000011101110011100101110 :
(key == 11'b01100111001) ? 46'b0001110110111010100101000011101101110101001010 :
(key == 11'b01100111010) ? 46'b0001110110100110110100000011101101001101101000 :
(key == 11'b01100111011) ? 46'b0001110110010011000100000011101100100110001000 :
(key == 11'b01100111100) ? 46'b0001110101111111010101000011101011111110101010 :
(key == 11'b01100111101) ? 46'b0001110101101011100111000011101011010111001110 :
(key == 11'b01100111110) ? 46'b0001110101010111111010000011101010101111110100 :
(key == 11'b01100111111) ? 46'b0001110101000100001110000011101010001000011100 :
(key == 11'b01101000000) ? 46'b0001110100110000100011000011101001100001000110 :
(key == 11'b01101000001) ? 46'b0001110100011100111001100011101000111001110011 :
(key == 11'b01101000010) ? 46'b0001110100001001010000100011101000010010100001 :
(key == 11'b01101000011) ? 46'b0001110011110101101000000011100111101011010000 :
(key == 11'b01101000100) ? 46'b0001110011100010000001100011100111000100000011 :
(key == 11'b01101000101) ? 46'b0001110011001110011011100011100110011100110111 :
(key == 11'b01101000110) ? 46'b0001110010111010110110100011100101110101101101 :
(key == 11'b01101000111) ? 46'b0001110010100111010011000011100101001110100110 :
(key == 11'b01101001000) ? 46'b0001110010010011110000000011100100100111100000 :
(key == 11'b01101001001) ? 46'b0001110010000000001110000011100100000000011100 :
(key == 11'b01101001010) ? 46'b0001110001101100101101000011100011011001011010 :
(key == 11'b01101001011) ? 46'b0001110001011001001101000011100010110010011010 :
(key == 11'b01101001100) ? 46'b0001110001000101101111000011100010001011011110 :
(key == 11'b01101001101) ? 46'b0001110000110010010001000011100001100100100010 :
(key == 11'b01101001110) ? 46'b0001110000011110110100000011100000111101101000 :
(key == 11'b01101001111) ? 46'b0001110000001011011000000011100000010110110000 :
(key == 11'b01101010000) ? 46'b0001101111110111111101000011011111101111111010 :
(key == 11'b01101010001) ? 46'b0001101111100100100011100011011111001001000111 :
(key == 11'b01101010010) ? 46'b0001101111010001001010100011011110100010010101 :
(key == 11'b01101010011) ? 46'b0001101110111101110011000011011101111011100110 :
(key == 11'b01101010100) ? 46'b0001101110101010011100000011011101010100111000 :
(key == 11'b01101010101) ? 46'b0001101110010111000110000011011100101110001100 :
(key == 11'b01101010110) ? 46'b0001101110000011110001000011011100000111100010 :
(key == 11'b01101010111) ? 46'b0001101101110000011101000011011011100000111010 :
(key == 11'b01101011000) ? 46'b0001101101011101001010000011011010111010010100 :
(key == 11'b01101011001) ? 46'b0001101101001001111000100011011010010011110001 :
(key == 11'b01101011010) ? 46'b0001101100110110100111100011011001101101001111 :
(key == 11'b01101011011) ? 46'b0001101100100011010111100011011001000110101111 :
(key == 11'b01101011100) ? 46'b0001101100010000001000100011011000100000010001 :
(key == 11'b01101011101) ? 46'b0001101011111100111010100011010111111001110101 :
(key == 11'b01101011110) ? 46'b0001101011101001101101100011010111010011011011 :
(key == 11'b01101011111) ? 46'b0001101011010110100001100011010110101101000011 :
(key == 11'b01101100000) ? 46'b0001101011000011010110100011010110000110101101 :
(key == 11'b01101100001) ? 46'b0001101010110000001100100011010101100000011001 :
(key == 11'b01101100010) ? 46'b0001101010011101000011100011010100111010000111 :
(key == 11'b01101100011) ? 46'b0001101010001001111011000011010100010011110110 :
(key == 11'b01101100100) ? 46'b0001101001110110110100000011010011101101101000 :
(key == 11'b01101100101) ? 46'b0001101001100011101110000011010011000111011100 :
(key == 11'b01101100110) ? 46'b0001101001010000101001000011010010100001010010 :
(key == 11'b01101100111) ? 46'b0001101000111101100100100011010001111011001001 :
(key == 11'b01101101000) ? 46'b0001101000101010100001000011010001010101000010 :
(key == 11'b01101101001) ? 46'b0001101000010111011111000011010000101110111110 :
(key == 11'b01101101010) ? 46'b0001101000000100011101100011010000001000111011 :
(key == 11'b01101101011) ? 46'b0001100111110001011100100011001111100010111001 :
(key == 11'b01101101100) ? 46'b0001100111011110011101000011001110111100111010 :
(key == 11'b01101101101) ? 46'b0001100111001011011111000011001110010110111110 :
(key == 11'b01101101110) ? 46'b0001100110111000100010000011001101110001000100 :
(key == 11'b01101101111) ? 46'b0001100110100101100101000011001101001011001010 :
(key == 11'b01101110000) ? 46'b0001100110010010101001000011001100100101010010 :
(key == 11'b01101110001) ? 46'b0001100101111111101110100011001011111111011101 :
(key == 11'b01101110010) ? 46'b0001100101101100110101000011001011011001101010 :
(key == 11'b01101110011) ? 46'b0001100101011001111100000011001010110011111000 :
(key == 11'b01101110100) ? 46'b0001100101000111000100000011001010001110001000 :
(key == 11'b01101110101) ? 46'b0001100100110100001101000011001001101000011010 :
(key == 11'b01101110110) ? 46'b0001100100100001010111000011001001000010101110 :
(key == 11'b01101110111) ? 46'b0001100100001110100010000011001000011101000100 :
(key == 11'b01101111000) ? 46'b0001100011111011101110100011000111110111011101 :
(key == 11'b01101111001) ? 46'b0001100011101000111011000011000111010001110110 :
(key == 11'b01101111010) ? 46'b0001100011010110001001000011000110101100010010 :
(key == 11'b01101111011) ? 46'b0001100011000011011000000011000110000110110000 :
(key == 11'b01101111100) ? 46'b0001100010110000101000000011000101100001010000 :
(key == 11'b01101111101) ? 46'b0001100010011101111000100011000100111011110001 :
(key == 11'b01101111110) ? 46'b0001100010001011001010000011000100010110010100 :
(key == 11'b01101111111) ? 46'b0001100001111000011100000011000011110000111000 :
(key == 11'b01110000000) ? 46'b0001100001100101110000000011000011001011100000 :
(key == 11'b01110000001) ? 46'b0001100001010011000100000011000010100110001000 :
(key == 11'b01110000010) ? 46'b0001100001000000011001100011000010000000110011 :
(key == 11'b01110000011) ? 46'b0001100000101101110000000011000001011011100000 :
(key == 11'b01110000100) ? 46'b0001100000011011000111000011000000110110001110 :
(key == 11'b01110000101) ? 46'b0001100000001000011111100011000000010000111111 :
(key == 11'b01110000110) ? 46'b0001011111110101111000100010111111101011110001 :
(key == 11'b01110000111) ? 46'b0001011111100011010010000010111111000110100100 :
(key == 11'b01110001000) ? 46'b0001011111010000101101000010111110100001011010 :
(key == 11'b01110001001) ? 46'b0001011110111110001001000010111101111100010010 :
(key == 11'b01110001010) ? 46'b0001011110101011100101100010111101010111001011 :
(key == 11'b01110001011) ? 46'b0001011110011001000011100010111100110010000111 :
(key == 11'b01110001100) ? 46'b0001011110000110100010000010111100001101000100 :
(key == 11'b01110001101) ? 46'b0001011101110100000010000010111011101000000100 :
(key == 11'b01110001110) ? 46'b0001011101100001100010000010111011000011000100 :
(key == 11'b01110001111) ? 46'b0001011101001111000011100010111010011110000111 :
(key == 11'b01110010000) ? 46'b0001011100111100100101100010111001111001001011 :
(key == 11'b01110010001) ? 46'b0001011100101010001001000010111001010100010010 :
(key == 11'b01110010010) ? 46'b0001011100010111101101000010111000101111011010 :
(key == 11'b01110010011) ? 46'b0001011100000101010010000010111000001010100100 :
(key == 11'b01110010100) ? 46'b0001011011110010111000000010110111100101110000 :
(key == 11'b01110010101) ? 46'b0001011011100000011111000010110111000000111110 :
(key == 11'b01110010110) ? 46'b0001011011001110000110100010110110011100001101 :
(key == 11'b01110010111) ? 46'b0001011010111011101111000010110101110111011110 :
(key == 11'b01110011000) ? 46'b0001011010101001011001000010110101010010110010 :
(key == 11'b01110011001) ? 46'b0001011010010111000011000010110100101110000110 :
(key == 11'b01110011010) ? 46'b0001011010000100101111000010110100001001011110 :
(key == 11'b01110011011) ? 46'b0001011001110010011011000010110011100100110110 :
(key == 11'b01110011100) ? 46'b0001011001100000001000000010110011000000010000 :
(key == 11'b01110011101) ? 46'b0001011001001101110110100010110010011011101101 :
(key == 11'b01110011110) ? 46'b0001011000111011100101000010110001110111001010 :
(key == 11'b01110011111) ? 46'b0001011000101001010101100010110001010010101011 :
(key == 11'b01110100000) ? 46'b0001011000010111000110000010110000101110001100 :
(key == 11'b01110100001) ? 46'b0001011000000100110111100010110000001001101111 :
(key == 11'b01110100010) ? 46'b0001010111110010101010000010101111100101010100 :
(key == 11'b01110100011) ? 46'b0001010111100000011101100010101111000000111011 :
(key == 11'b01110100100) ? 46'b0001010111001110010010000010101110011100100100 :
(key == 11'b01110100101) ? 46'b0001010110111100000111000010101101111000001110 :
(key == 11'b01110100110) ? 46'b0001010110101001111101000010101101010011111010 :
(key == 11'b01110100111) ? 46'b0001010110010111110100000010101100101111101000 :
(key == 11'b01110101000) ? 46'b0001010110000101101100000010101100001011011000 :
(key == 11'b01110101001) ? 46'b0001010101110011100101000010101011100111001010 :
(key == 11'b01110101010) ? 46'b0001010101100001011111000010101011000010111110 :
(key == 11'b01110101011) ? 46'b0001010101001111011010000010101010011110110100 :
(key == 11'b01110101100) ? 46'b0001010100111101010101000010101001111010101010 :
(key == 11'b01110101101) ? 46'b0001010100101011010001100010101001010110100011 :
(key == 11'b01110101110) ? 46'b0001010100011001001110100010101000110010011101 :
(key == 11'b01110101111) ? 46'b0001010100000111001100100010101000001110011001 :
(key == 11'b01110110000) ? 46'b0001010011110101001011100010100111101010010111 :
(key == 11'b01110110001) ? 46'b0001010011100011001011100010100111000110010111 :
(key == 11'b01110110010) ? 46'b0001010011010001001100000010100110100010011000 :
(key == 11'b01110110011) ? 46'b0001010010111111001110000010100101111110011100 :
(key == 11'b01110110100) ? 46'b0001010010101101010000100010100101011010100001 :
(key == 11'b01110110101) ? 46'b0001010010011011010100000010100100110110101000 :
(key == 11'b01110110110) ? 46'b0001010010001001011000000010100100010010110000 :
(key == 11'b01110110111) ? 46'b0001010001110111011101000010100011101110111010 :
(key == 11'b01110111000) ? 46'b0001010001100101100011000010100011001011000110 :
(key == 11'b01110111001) ? 46'b0001010001010011101010000010100010100111010100 :
(key == 11'b01110111010) ? 46'b0001010001000001110010000010100010000011100100 :
(key == 11'b01110111011) ? 46'b0001010000101111111010000010100001011111110100 :
(key == 11'b01110111100) ? 46'b0001010000011110000100000010100000111100001000 :
(key == 11'b01110111101) ? 46'b0001010000001100001110000010100000011000011100 :
(key == 11'b01110111110) ? 46'b0001001111111010011001100010011111110100110011 :
(key == 11'b01110111111) ? 46'b0001001111101000100101100010011111010001001011 :
(key == 11'b01111000000) ? 46'b0001001111010110110010000010011110101101100100 :
(key == 11'b01111000001) ? 46'b0001001111000101000000000010011110001010000000 :
(key == 11'b01111000010) ? 46'b0001001110110011001110100010011101100110011101 :
(key == 11'b01111000011) ? 46'b0001001110100001011110000010011101000010111100 :
(key == 11'b01111000100) ? 46'b0001001110001111101110000010011100011111011100 :
(key == 11'b01111000101) ? 46'b0001001101111101111111100010011011111011111111 :
(key == 11'b01111000110) ? 46'b0001001101101100010001100010011011011000100011 :
(key == 11'b01111000111) ? 46'b0001001101011010100100000010011010110101001000 :
(key == 11'b01111001000) ? 46'b0001001101001000111000000010011010010001110000 :
(key == 11'b01111001001) ? 46'b0001001100110111001101000010011001101110011010 :
(key == 11'b01111001010) ? 46'b0001001100100101100010000010011001001011000100 :
(key == 11'b01111001011) ? 46'b0001001100010011111000000010011000100111110000 :
(key == 11'b01111001100) ? 46'b0001001100000010001111100010011000000100011111 :
(key == 11'b01111001101) ? 46'b0001001011110000100111100010010111100001001111 :
(key == 11'b01111001110) ? 46'b0001001011011111000000100010010110111110000001 :
(key == 11'b01111001111) ? 46'b0001001011001101011010100010010110011010110101 :
(key == 11'b01111010000) ? 46'b0001001010111011110101000010010101110111101010 :
(key == 11'b01111010001) ? 46'b0001001010101010010000100010010101010100100001 :
(key == 11'b01111010010) ? 46'b0001001010011000101100100010010100110001011001 :
(key == 11'b01111010011) ? 46'b0001001010000111001001100010010100001110010011 :
(key == 11'b01111010100) ? 46'b0001001001110101100111100010010011101011001111 :
(key == 11'b01111010101) ? 46'b0001001001100100000110000010010011001000001100 :
(key == 11'b01111010110) ? 46'b0001001001010010100110000010010010100101001100 :
(key == 11'b01111010111) ? 46'b0001001001000001000110000010010010000010001100 :
(key == 11'b01111011000) ? 46'b0001001000101111101000000010010001011111010000 :
(key == 11'b01111011001) ? 46'b0001001000011110001010000010010000111100010100 :
(key == 11'b01111011010) ? 46'b0001001000001100101101000010010000011001011010 :
(key == 11'b01111011011) ? 46'b0001000111111011010000100010001111110110100001 :
(key == 11'b01111011100) ? 46'b0001000111101001110101000010001111010011101010 :
(key == 11'b01111011101) ? 46'b0001000111011000011010000010001110110000110100 :
(key == 11'b01111011110) ? 46'b0001000111000111000000100010001110001110000001 :
(key == 11'b01111011111) ? 46'b0001000110110101101000000010001101101011010000 :
(key == 11'b01111100000) ? 46'b0001000110100100010000000010001101001000100000 :
(key == 11'b01111100001) ? 46'b0001000110010010111000100010001100100101110001 :
(key == 11'b01111100010) ? 46'b0001000110000001100010000010001100000011000100 :
(key == 11'b01111100011) ? 46'b0001000101110000001100100010001011100000011001 :
(key == 11'b01111100100) ? 46'b0001000101011110111000000010001010111101110000 :
(key == 11'b01111100101) ? 46'b0001000101001101100100000010001010011011001000 :
(key == 11'b01111100110) ? 46'b0001000100111100010000100010001001111000100001 :
(key == 11'b01111100111) ? 46'b0001000100101010111110000010001001010101111100 :
(key == 11'b01111101000) ? 46'b0001000100011001101101000010001000110011011010 :
(key == 11'b01111101001) ? 46'b0001000100001000011100000010001000010000111000 :
(key == 11'b01111101010) ? 46'b0001000011110111001100000010000111101110011000 :
(key == 11'b01111101011) ? 46'b0001000011100101111101000010000111001011111010 :
(key == 11'b01111101100) ? 46'b0001000011010100101111000010000110101001011110 :
(key == 11'b01111101101) ? 46'b0001000011000011100001100010000110000111000011 :
(key == 11'b01111101110) ? 46'b0001000010110010010101000010000101100100101010 :
(key == 11'b01111101111) ? 46'b0001000010100001001001100010000101000010010011 :
(key == 11'b01111110000) ? 46'b0001000010001111111110100010000100011111111101 :
(key == 11'b01111110001) ? 46'b0001000001111110110100000010000011111101101000 :
(key == 11'b01111110010) ? 46'b0001000001101101101011000010000011011011010110 :
(key == 11'b01111110011) ? 46'b0001000001011100100010000010000010111001000100 :
(key == 11'b01111110100) ? 46'b0001000001001011011010100010000010010110110101 :
(key == 11'b01111110101) ? 46'b0001000000111010010011100010000001110100100111 :
(key == 11'b01111110110) ? 46'b0001000000101001001101000010000001010010011010 :
(key == 11'b01111110111) ? 46'b0001000000011000001000000010000000110000010000 :
(key == 11'b01111111000) ? 46'b0001000000000111000100000010000000001110001000 :
(key == 11'b01111111001) ? 46'b0000111111110110000000000001111111101100000000 :
(key == 11'b01111111010) ? 46'b0000111111100100111101000001111111001001111010 :
(key == 11'b01111111011) ? 46'b0000111111010011111011000001111110100111110110 :
(key == 11'b01111111100) ? 46'b0000111111000010111010000001111110000101110100 :
(key == 11'b01111111101) ? 46'b0000111110110001111001000001111101100011110010 :
(key == 11'b01111111110) ? 46'b0000111110100000111001000001111101000001110010 :
(key == 11'b01111111111) ? 46'b0000111110001111111010100001111100011111110101 :
(key == 11'b10000000000) ? 46'b0111111111101000000001001111111111010000000010 :
(key == 11'b10000000001) ? 46'b0111111110111000000101101111111101110000001011 :
(key == 11'b10000000010) ? 46'b0111111110001000001111001111111100010000011110 :
(key == 11'b10000000011) ? 46'b0111111101011000011100001111111010110000111000 :
(key == 11'b10000000100) ? 46'b0111111100101000101110001111111001010001011100 :
(key == 11'b10000000101) ? 46'b0111111011111001000100101111110111110010001001 :
(key == 11'b10000000110) ? 46'b0111111011001001011111101111110110010010111111 :
(key == 11'b10000000111) ? 46'b0111111010011001111110101111110100110011111101 :
(key == 11'b10000001000) ? 46'b0111111001101010100010101111110011010101000101 :
(key == 11'b10000001001) ? 46'b0111111000111011001010001111110001110110010100 :
(key == 11'b10000001010) ? 46'b0111111000001011110111001111110000010111101110 :
(key == 11'b10000001011) ? 46'b0111110111011100100111101111101110111001001111 :
(key == 11'b10000001100) ? 46'b0111110110101101011100101111101101011010111001 :
(key == 11'b10000001101) ? 46'b0111110101111110010110001111101011111100101100 :
(key == 11'b10000001110) ? 46'b0111110101001111010011101111101010011110100111 :
(key == 11'b10000001111) ? 46'b0111110100100000010110101111101001000000101101 :
(key == 11'b10000010000) ? 46'b0111110011110001011101001111100111100010111010 :
(key == 11'b10000010001) ? 46'b0111110011000010101000001111100110000101010000 :
(key == 11'b10000010010) ? 46'b0111110010010011111000001111100100100111110000 :
(key == 11'b10000010011) ? 46'b0111110001100101001010101111100011001010010101 :
(key == 11'b10000010100) ? 46'b0111110000110110100011001111100001101101000110 :
(key == 11'b10000010101) ? 46'b0111110000000111111110101111100000001111111101 :
(key == 11'b10000010110) ? 46'b0111101111011001011111101111011110110010111111 :
(key == 11'b10000010111) ? 46'b0111101110101011000011101111011101010110000111 :
(key == 11'b10000011000) ? 46'b0111101101111100101101001111011011111001011010 :
(key == 11'b10000011001) ? 46'b0111101101001110011010101111011010011100110101 :
(key == 11'b10000011010) ? 46'b0111101100100000001011001111011001000000010110 :
(key == 11'b10000011011) ? 46'b0111101011110010000001101111010111100100000011 :
(key == 11'b10000011100) ? 46'b0111101011000011111010101111010110000111110101 :
(key == 11'b10000011101) ? 46'b0111101010010101111001001111010100101011110010 :
(key == 11'b10000011110) ? 46'b0111101001100111111010101111010011001111110101 :
(key == 11'b10000011111) ? 46'b0111101000111010000001101111010001110100000011 :
(key == 11'b10000100000) ? 46'b0111101000001100001100001111010000011000011000 :
(key == 11'b10000100001) ? 46'b0111100111011110011010101111001110111100110101 :
(key == 11'b10000100010) ? 46'b0111100110110000101110001111001101100001011100 :
(key == 11'b10000100011) ? 46'b0111100110000011000100101111001100000110001001 :
(key == 11'b10000100100) ? 46'b0111100101010101100000001111001010101011000000 :
(key == 11'b10000100101) ? 46'b0111100100100111111111001111001001001111111110 :
(key == 11'b10000100110) ? 46'b0111100011111010100010101111000111110101000101 :
(key == 11'b10000100111) ? 46'b0111100011001101001010101111000110011010010101 :
(key == 11'b10000101000) ? 46'b0111100010011111110101101111000100111111101011 :
(key == 11'b10000101001) ? 46'b0111100001110010100101101111000011100101001011 :
(key == 11'b10000101010) ? 46'b0111100001000101011001001111000010001010110010 :
(key == 11'b10000101011) ? 46'b0111100000011000010001101111000000110000100011 :
(key == 11'b10000101100) ? 46'b0111011111101011001100001110111111010110011000 :
(key == 11'b10000101101) ? 46'b0111011110111110001100101110111101111100011001 :
(key == 11'b10000101110) ? 46'b0111011110010001010000001110111100100010100000 :
(key == 11'b10000101111) ? 46'b0111011101100100011001001110111011001000110010 :
(key == 11'b10000110000) ? 46'b0111011100110111100101001110111001101111001010 :
(key == 11'b10000110001) ? 46'b0111011100001010110100101110111000010101101001 :
(key == 11'b10000110010) ? 46'b0111011011011110001000101110110110111100010001 :
(key == 11'b10000110011) ? 46'b0111011010110001100001001110110101100011000010 :
(key == 11'b10000110100) ? 46'b0111011010000100111101001110110100001001111010 :
(key == 11'b10000110101) ? 46'b0111011001011000011100101110110010110000111001 :
(key == 11'b10000110110) ? 46'b0111011000101100000000101110110001011000000001 :
(key == 11'b10000110111) ? 46'b0111010111111111101000101110101111111111010001 :
(key == 11'b10000111000) ? 46'b0111010111010011010100001110101110100110101000 :
(key == 11'b10000111001) ? 46'b0111010110100111000100001110101101001110001000 :
(key == 11'b10000111010) ? 46'b0111010101111010110111001110101011110101101110 :
(key == 11'b10000111011) ? 46'b0111010101001110101111001110101010011101011110 :
(key == 11'b10000111100) ? 46'b0111010100100010101010001110101001000101010100 :
(key == 11'b10000111101) ? 46'b0111010011110110101010001110100111101101010100 :
(key == 11'b10000111110) ? 46'b0111010011001010101101001110100110010101011010 :
(key == 11'b10000111111) ? 46'b0111010010011110110101001110100100111101101010 :
(key == 11'b10001000000) ? 46'b0111010001110011000000001110100011100110000000 :
(key == 11'b10001000001) ? 46'b0111010001000111001110001110100010001110011100 :
(key == 11'b10001000010) ? 46'b0111010000011011100001001110100000110111000010 :
(key == 11'b10001000011) ? 46'b0111001111101111110111101110011111011111101111 :
(key == 11'b10001000100) ? 46'b0111001111000100010001101110011110001000100011 :
(key == 11'b10001000101) ? 46'b0111001110011000110000101110011100110001100001 :
(key == 11'b10001000110) ? 46'b0111001101101101010010101110011011011010100101 :
(key == 11'b10001000111) ? 46'b0111001101000001111000101110011010000011110001 :
(key == 11'b10001001000) ? 46'b0111001100010110100010001110011000101101000100 :
(key == 11'b10001001001) ? 46'b0111001011101011001111001110010111010110011110 :
(key == 11'b10001001010) ? 46'b0111001011000000000001001110010110000000000010 :
(key == 11'b10001001011) ? 46'b0111001010010100110110001110010100101001101100 :
(key == 11'b10001001100) ? 46'b0111001001101001101110101110010011010011011101 :
(key == 11'b10001001101) ? 46'b0111001000111110101011001110010001111101010110 :
(key == 11'b10001001110) ? 46'b0111001000010011101011101110010000100111010111 :
(key == 11'b10001001111) ? 46'b0111000111101000110000001110001111010001100000 :
(key == 11'b10001010000) ? 46'b0111000110111101110111001110001101111011101110 :
(key == 11'b10001010001) ? 46'b0111000110010011000011001110001100100110000110 :
(key == 11'b10001010010) ? 46'b0111000101101000010010001110001011010000100100 :
(key == 11'b10001010011) ? 46'b0111000100111101100101001110001001111011001010 :
(key == 11'b10001010100) ? 46'b0111000100010010111011101110001000100101110111 :
(key == 11'b10001010101) ? 46'b0111000011101000010110001110000111010000101100 :
(key == 11'b10001010110) ? 46'b0111000010111101110100001110000101111011101000 :
(key == 11'b10001010111) ? 46'b0111000010010011010101101110000100100110101011 :
(key == 11'b10001011000) ? 46'b0111000001101000111011101110000011010001110111 :
(key == 11'b10001011001) ? 46'b0111000000111110100100001110000001111101001000 :
(key == 11'b10001011010) ? 46'b0111000000010100010000001110000000101000100000 :
(key == 11'b10001011011) ? 46'b0110111111101010000001001101111111010100000010 :
(key == 11'b10001011100) ? 46'b0110111110111111110101001101111101111111101010 :
(key == 11'b10001011101) ? 46'b0110111110010101101100001101111100101011011000 :
(key == 11'b10001011110) ? 46'b0110111101101011100111001101111011010111001110 :
(key == 11'b10001011111) ? 46'b0110111101000001100110001101111010000011001100 :
(key == 11'b10001100000) ? 46'b0110111100010111101001001101111000101111010010 :
(key == 11'b10001100001) ? 46'b0110111011101101101111001101110111011011011110 :
(key == 11'b10001100010) ? 46'b0110111011000011111000001101110110000111110000 :
(key == 11'b10001100011) ? 46'b0110111010011010000101001101110100110100001010 :
(key == 11'b10001100100) ? 46'b0110111001110000010110001101110011100000101100 :
(key == 11'b10001100101) ? 46'b0110111001000110101010101101110010001101010101 :
(key == 11'b10001100110) ? 46'b0110111000011101000010101101110000111010000101 :
(key == 11'b10001100111) ? 46'b0110110111110011011101001101101111100110111010 :
(key == 11'b10001101000) ? 46'b0110110111001001111100001101101110010011111000 :
(key == 11'b10001101001) ? 46'b0110110110100000011111001101101101000000111110 :
(key == 11'b10001101010) ? 46'b0110110101110111000101001101101011101110001010 :
(key == 11'b10001101011) ? 46'b0110110101001101101110001101101010011011011100 :
(key == 11'b10001101100) ? 46'b0110110100100100011011101101101001001000110111 :
(key == 11'b10001101101) ? 46'b0110110011111011001011101101100111110110010111 :
(key == 11'b10001101110) ? 46'b0110110011010010000000001101100110100100000000 :
(key == 11'b10001101111) ? 46'b0110110010101000110111001101100101010001101110 :
(key == 11'b10001110000) ? 46'b0110110001111111110010001101100011111111100100 :
(key == 11'b10001110001) ? 46'b0110110001010110110000101101100010101101100001 :
(key == 11'b10001110010) ? 46'b0110110000101101110010101101100001011011100101 :
(key == 11'b10001110011) ? 46'b0110110000000100111000001101100000001001110000 :
(key == 11'b10001110100) ? 46'b0110101111011100000000101101011110111000000001 :
(key == 11'b10001110101) ? 46'b0110101110110011001100101101011101100110011001 :
(key == 11'b10001110110) ? 46'b0110101110001010011100001101011100010100111000 :
(key == 11'b10001110111) ? 46'b0110101101100001101111001101011011000011011110 :
(key == 11'b10001111000) ? 46'b0110101100111001000101101101011001110010001011 :
(key == 11'b10001111001) ? 46'b0110101100010000011111101101011000100000111111 :
(key == 11'b10001111010) ? 46'b0110101011100111111100101101010111001111111001 :
(key == 11'b10001111011) ? 46'b0110101010111111011101001101010101111110111010 :
(key == 11'b10001111100) ? 46'b0110101010010111000001101101010100101110000011 :
(key == 11'b10001111101) ? 46'b0110101001101110101001001101010011011101010010 :
(key == 11'b10001111110) ? 46'b0110101001000110010011101101010010001100100111 :
(key == 11'b10001111111) ? 46'b0110101000011110000010001101010000111100000100 :
(key == 11'b10010000000) ? 46'b0110100111110101110011101101001111101011100111 :
(key == 11'b10010000001) ? 46'b0110100111001101100111101101001110011011001111 :
(key == 11'b10010000010) ? 46'b0110100110100101100000101101001101001011000001 :
(key == 11'b10010000011) ? 46'b0110100101111101011100001101001011111010111000 :
(key == 11'b10010000100) ? 46'b0110100101010101011011001101001010101010110110 :
(key == 11'b10010000101) ? 46'b0110100100101101011101001101001001011010111010 :
(key == 11'b10010000110) ? 46'b0110100100000101100010101101001000001011000101 :
(key == 11'b10010000111) ? 46'b0110100011011101101011101101000110111011010111 :
(key == 11'b10010001000) ? 46'b0110100010110101110111101101000101101011101111 :
(key == 11'b10010001001) ? 46'b0110100010001110000111001101000100011100001110 :
(key == 11'b10010001010) ? 46'b0110100001100110011001101101000011001100110011 :
(key == 11'b10010001011) ? 46'b0110100000111110101111001101000001111101011110 :
(key == 11'b10010001100) ? 46'b0110100000010111001001001101000000101110010010 :
(key == 11'b10010001101) ? 46'b0110011111101111100101001100111111011111001010 :
(key == 11'b10010001110) ? 46'b0110011111001000000100001100111110010000001000 :
(key == 11'b10010001111) ? 46'b0110011110100000100111101100111101000001001111 :
(key == 11'b10010010000) ? 46'b0110011101111001001110001100111011110010011100 :
(key == 11'b10010010001) ? 46'b0110011101010001110111101100111010100011101111 :
(key == 11'b10010010010) ? 46'b0110011100101010100100001100111001010101001000 :
(key == 11'b10010010011) ? 46'b0110011100000011010100001100111000000110101000 :
(key == 11'b10010010100) ? 46'b0110011011011100000110101100110110111000001101 :
(key == 11'b10010010101) ? 46'b0110011010110100111101001100110101101001111010 :
(key == 11'b10010010110) ? 46'b0110011010001101110111001100110100011011101110 :
(key == 11'b10010010111) ? 46'b0110011001100110110011101100110011001101100111 :
(key == 11'b10010011000) ? 46'b0110011000111111110011101100110001111111100111 :
(key == 11'b10010011001) ? 46'b0110011000011000110111001100110000110001101110 :
(key == 11'b10010011010) ? 46'b0110010111110001111101001100101111100011111010 :
(key == 11'b10010011011) ? 46'b0110010111001011000110001100101110010110001100 :
(key == 11'b10010011100) ? 46'b0110010110100100010011001100101101001000100110 :
(key == 11'b10010011101) ? 46'b0110010101111101100010101100101011111011000101 :
(key == 11'b10010011110) ? 46'b0110010101010110110110001100101010101101101100 :
(key == 11'b10010011111) ? 46'b0110010100110000001011001100101001100000010110 :
(key == 11'b10010100000) ? 46'b0110010100001001100101001100101000010011001010 :
(key == 11'b10010100001) ? 46'b0110010011100011000001001100100111000110000010 :
(key == 11'b10010100010) ? 46'b0110010010111100100000101100100101111001000001 :
(key == 11'b10010100011) ? 46'b0110010010010110000011001100100100101100000110 :
(key == 11'b10010100100) ? 46'b0110010001101111101001001100100011011111010010 :
(key == 11'b10010100101) ? 46'b0110010001001001010001001100100010010010100010 :
(key == 11'b10010100110) ? 46'b0110010000100010111101001100100001000101111010 :
(key == 11'b10010100111) ? 46'b0110001111111100101100001100011111111001011000 :
(key == 11'b10010101000) ? 46'b0110001111010110011110001100011110101100111100 :
(key == 11'b10010101001) ? 46'b0110001110110000010011101100011101100000100111 :
(key == 11'b10010101010) ? 46'b0110001110001010001011101100011100010100010111 :
(key == 11'b10010101011) ? 46'b0110001101100100000110001100011011001000001100 :
(key == 11'b10010101100) ? 46'b0110001100111110000101001100011001111100001010 :
(key == 11'b10010101101) ? 46'b0110001100011000000110001100011000110000001100 :
(key == 11'b10010101110) ? 46'b0110001011110010001010101100010111100100010101 :
(key == 11'b10010101111) ? 46'b0110001011001100010001101100010110011000100011 :
(key == 11'b10010110000) ? 46'b0110001010100110011100001100010101001100111000 :
(key == 11'b10010110001) ? 46'b0110001010000000101010001100010100000001010100 :
(key == 11'b10010110010) ? 46'b0110001001011010111010001100010010110101110100 :
(key == 11'b10010110011) ? 46'b0110001000110101001101101100010001101010011011 :
(key == 11'b10010110100) ? 46'b0110001000001111100100001100010000011111001000 :
(key == 11'b10010110101) ? 46'b0110000111101001111101001100001111010011111010 :
(key == 11'b10010110110) ? 46'b0110000111000100011010001100001110001000110100 :
(key == 11'b10010110111) ? 46'b0110000110011110111001101100001100111101110011 :
(key == 11'b10010111000) ? 46'b0110000101111001011011101100001011110010110111 :
(key == 11'b10010111001) ? 46'b0110000101010100000001001100001010101000000010 :
(key == 11'b10010111010) ? 46'b0110000100101110101001101100001001011101010011 :
(key == 11'b10010111011) ? 46'b0110000100001001010101001100001000010010101010 :
(key == 11'b10010111100) ? 46'b0110000011100100000011001100000111001000000110 :
(key == 11'b10010111101) ? 46'b0110000010111110110100101100000101111101101001 :
(key == 11'b10010111110) ? 46'b0110000010011001101000101100000100110011010001 :
(key == 11'b10010111111) ? 46'b0110000001110100100000001100000011101001000000 :
(key == 11'b10011000000) ? 46'b0110000001001111011010001100000010011110110100 :
(key == 11'b10011000001) ? 46'b0110000000101010010111001100000001010100101110 :
(key == 11'b10011000010) ? 46'b0110000000000101010110101100000000001010101101 :
(key == 11'b10011000011) ? 46'b0101111111100000011001101011111111000000110011 :
(key == 11'b10011000100) ? 46'b0101111110111011011111001011111101110110111110 :
(key == 11'b10011000101) ? 46'b0101111110010110101000001011111100101101010000 :
(key == 11'b10011000110) ? 46'b0101111101110001110011101011111011100011100111 :
(key == 11'b10011000111) ? 46'b0101111101001101000010001011111010011010000100 :
(key == 11'b10011001000) ? 46'b0101111100101000010011001011111001010000100110 :
(key == 11'b10011001001) ? 46'b0101111100000011100111001011111000000111001110 :
(key == 11'b10011001010) ? 46'b0101111011011110111110001011110110111101111100 :
(key == 11'b10011001011) ? 46'b0101111010111010011000001011110101110100110000 :
(key == 11'b10011001100) ? 46'b0101111010010101110101001011110100101011101010 :
(key == 11'b10011001101) ? 46'b0101111001110001010101001011110011100010101010 :
(key == 11'b10011001110) ? 46'b0101111001001100110111001011110010011001101110 :
(key == 11'b10011001111) ? 46'b0101111000101000011100101011110001010000111001 :
(key == 11'b10011010000) ? 46'b0101111000000100000101001011110000001000001010 :
(key == 11'b10011010001) ? 46'b0101110111011111101111101011101110111111011111 :
(key == 11'b10011010010) ? 46'b0101110110111011011101001011101101110110111010 :
(key == 11'b10011010011) ? 46'b0101110110010111001110101011101100101110011101 :
(key == 11'b10011010100) ? 46'b0101110101110011000001101011101011100110000011 :
(key == 11'b10011010101) ? 46'b0101110101001110110111101011101010011101101111 :
(key == 11'b10011010110) ? 46'b0101110100101010110000101011101001010101100001 :
(key == 11'b10011010111) ? 46'b0101110100000110101100101011101000001101011001 :
(key == 11'b10011011000) ? 46'b0101110011100010101011001011100111000101010110 :
(key == 11'b10011011001) ? 46'b0101110010111110101100101011100101111101011001 :
(key == 11'b10011011010) ? 46'b0101110010011010110000101011100100110101100001 :
(key == 11'b10011011011) ? 46'b0101110001110110111000001011100011101101110000 :
(key == 11'b10011011100) ? 46'b0101110001010011000010001011100010100110000100 :
(key == 11'b10011011101) ? 46'b0101110000101111001110001011100001011110011100 :
(key == 11'b10011011110) ? 46'b0101110000001011011101001011100000010110111010 :
(key == 11'b10011011111) ? 46'b0101101111100111101111001011011111001111011110 :
(key == 11'b10011100000) ? 46'b0101101111000100000100101011011110001000001001 :
(key == 11'b10011100001) ? 46'b0101101110100000011100001011011101000000111000 :
(key == 11'b10011100010) ? 46'b0101101101111100110110001011011011111001101100 :
(key == 11'b10011100011) ? 46'b0101101101011001010011001011011010110010100110 :
(key == 11'b10011100100) ? 46'b0101101100110101110011001011011001101011100110 :
(key == 11'b10011100101) ? 46'b0101101100010010010101001011011000100100101010 :
(key == 11'b10011100110) ? 46'b0101101011101110111010101011010111011101110101 :
(key == 11'b10011100111) ? 46'b0101101011001011100010001011010110010111000100 :
(key == 11'b10011101000) ? 46'b0101101010101000001100101011010101010000011001 :
(key == 11'b10011101001) ? 46'b0101101010000100111010001011010100001001110100 :
(key == 11'b10011101010) ? 46'b0101101001100001101010001011010011000011010100 :
(key == 11'b10011101011) ? 46'b0101101000111110011100101011010001111100111001 :
(key == 11'b10011101100) ? 46'b0101101000011011010010001011010000110110100100 :
(key == 11'b10011101101) ? 46'b0101100111111000001001101011001111110000010011 :
(key == 11'b10011101110) ? 46'b0101100111010101000101001011001110101010001010 :
(key == 11'b10011101111) ? 46'b0101100110110010000001101011001101100100000011 :
(key == 11'b10011110000) ? 46'b0101100110001111000001101011001100011110000011 :
(key == 11'b10011110001) ? 46'b0101100101101100000100101011001011011000001001 :
(key == 11'b10011110010) ? 46'b0101100101001001001001101011001010010010010011 :
(key == 11'b10011110011) ? 46'b0101100100100110010001001011001001001100100010 :
(key == 11'b10011110100) ? 46'b0101100100000011011100001011001000000110111000 :
(key == 11'b10011110101) ? 46'b0101100011100000101010001011000111000001010100 :
(key == 11'b10011110110) ? 46'b0101100010111101111001001011000101111011110010 :
(key == 11'b10011110111) ? 46'b0101100010011011001100001011000100110110011000 :
(key == 11'b10011111000) ? 46'b0101100001111000100000101011000011110001000001 :
(key == 11'b10011111001) ? 46'b0101100001010101111000001011000010101011110000 :
(key == 11'b10011111010) ? 46'b0101100000110011010010101011000001100110100101 :
(key == 11'b10011111011) ? 46'b0101100000010000101111101011000000100001011111 :
(key == 11'b10011111100) ? 46'b0101011111101110001111001010111111011100011110 :
(key == 11'b10011111101) ? 46'b0101011111001011110001001010111110010111100010 :
(key == 11'b10011111110) ? 46'b0101011110101001010101101010111101010010101011 :
(key == 11'b10011111111) ? 46'b0101011110000110111101001010111100001101111010 :
(key == 11'b10100000000) ? 46'b0101011101100100100111001010111011001001001110 :
(key == 11'b10100000001) ? 46'b0101011101000010010011101010111010000100100111 :
(key == 11'b10100000010) ? 46'b0101011100100000000010001010111001000000000100 :
(key == 11'b10100000011) ? 46'b0101011011111101110100001010110111111011101000 :
(key == 11'b10100000100) ? 46'b0101011011011011101000001010110110110111010000 :
(key == 11'b10100000101) ? 46'b0101011010111001011110101010110101110010111101 :
(key == 11'b10100000110) ? 46'b0101011010010111011000001010110100101110110000 :
(key == 11'b10100000111) ? 46'b0101011001110101010011101010110011101010100111 :
(key == 11'b10100001000) ? 46'b0101011001010011010010001010110010100110100100 :
(key == 11'b10100001001) ? 46'b0101011000110001010011001010110001100010100110 :
(key == 11'b10100001010) ? 46'b0101011000001111010110001010110000011110101100 :
(key == 11'b10100001011) ? 46'b0101010111101101011100001010101111011010111000 :
(key == 11'b10100001100) ? 46'b0101010111001011100101001010101110010111001010 :
(key == 11'b10100001101) ? 46'b0101010110101001101111001010101101010011011110 :
(key == 11'b10100001110) ? 46'b0101010110000111111100001010101100001111111000 :
(key == 11'b10100001111) ? 46'b0101010101100110001101001010101011001100011010 :
(key == 11'b10100010000) ? 46'b0101010101000100011111001010101010001000111110 :
(key == 11'b10100010001) ? 46'b0101010100100010110100001010101001000101101000 :
(key == 11'b10100010010) ? 46'b0101010100000001001011001010101000000010010110 :
(key == 11'b10100010011) ? 46'b0101010011011111100101001010100110111111001010 :
(key == 11'b10100010100) ? 46'b0101010010111110000010001010100101111100000100 :
(key == 11'b10100010101) ? 46'b0101010010011100100001001010100100111001000010 :
(key == 11'b10100010110) ? 46'b0101010001111011000010001010100011110110000100 :
(key == 11'b10100010111) ? 46'b0101010001011001100101101010100010110011001011 :
(key == 11'b10100011000) ? 46'b0101010000111000001100101010100001110000011001 :
(key == 11'b10100011001) ? 46'b0101010000010110110101001010100000101101101010 :
(key == 11'b10100011010) ? 46'b0101001111110101100000101010011111101011000001 :
(key == 11'b10100011011) ? 46'b0101001111010100001101101010011110101000011011 :
(key == 11'b10100011100) ? 46'b0101001110110010111101101010011101100101111011 :
(key == 11'b10100011101) ? 46'b0101001110010001110000001010011100100011100000 :
(key == 11'b10100011110) ? 46'b0101001101110000100101001010011011100001001010 :
(key == 11'b10100011111) ? 46'b0101001101001111011100101010011010011110111001 :
(key == 11'b10100100000) ? 46'b0101001100101110010110001010011001011100101100 :
(key == 11'b10100100001) ? 46'b0101001100001101010010101010011000011010100101 :
(key == 11'b10100100010) ? 46'b0101001011101100010001001010010111011000100010 :
(key == 11'b10100100011) ? 46'b0101001011001011010010001010010110010110100100 :
(key == 11'b10100100100) ? 46'b0101001010101010010110001010010101010100101100 :
(key == 11'b10100100101) ? 46'b0101001010001001011100001010010100010010111000 :
(key == 11'b10100100110) ? 46'b0101001001101000100011101010010011010001000111 :
(key == 11'b10100100111) ? 46'b0101001001000111101110001010010010001111011100 :
(key == 11'b10100101000) ? 46'b0101001000100110111011101010010001001101110111 :
(key == 11'b10100101001) ? 46'b0101001000000110001010101010010000001100010101 :
(key == 11'b10100101010) ? 46'b0101000111100101011100101010001111001010111001 :
(key == 11'b10100101011) ? 46'b0101000111000100110000001010001110001001100000 :
(key == 11'b10100101100) ? 46'b0101000110100100000111101010001101001000001111 :
(key == 11'b10100101101) ? 46'b0101000110000011100000001010001100000111000000 :
(key == 11'b10100101110) ? 46'b0101000101100010111011001010001011000101110110 :
(key == 11'b10100101111) ? 46'b0101000101000010011001001010001010000100110010 :
(key == 11'b10100110000) ? 46'b0101000100100001111001001010001001000011110010 :
(key == 11'b10100110001) ? 46'b0101000100000001011011001010001000000010110110 :
(key == 11'b10100110010) ? 46'b0101000011100000111111101010000111000001111111 :
(key == 11'b10100110011) ? 46'b0101000011000000100110101010000110000001001101 :
(key == 11'b10100110100) ? 46'b0101000010100000010000001010000101000000100000 :
(key == 11'b10100110101) ? 46'b0101000001111111111011101010000011111111110111 :
(key == 11'b10100110110) ? 46'b0101000001011111101010001010000010111111010100 :
(key == 11'b10100110111) ? 46'b0101000000111111011010001010000001111110110100 :
(key == 11'b10100111000) ? 46'b0101000000011111001101001010000000111110011010 :
(key == 11'b10100111001) ? 46'b0100111111111111000001001001111111111110000010 :
(key == 11'b10100111010) ? 46'b0100111111011110111000101001111110111101110001 :
(key == 11'b10100111011) ? 46'b0100111110111110110010001001111101111101100100 :
(key == 11'b10100111100) ? 46'b0100111110011110101110001001111100111101011100 :
(key == 11'b10100111101) ? 46'b0100111101111110101100101001111011111101011001 :
(key == 11'b10100111110) ? 46'b0100111101011110101100001001111010111101011000 :
(key == 11'b10100111111) ? 46'b0100111100111110101111101001111001111101011111 :
(key == 11'b10101000000) ? 46'b0100111100011110110100101001111000111101101001 :
(key == 11'b10101000001) ? 46'b0100111011111110111011001001110111111101110110 :
(key == 11'b10101000010) ? 46'b0100111011011111000101001001110110111110001010 :
(key == 11'b10101000011) ? 46'b0100111010111111010001001001110101111110100010 :
(key == 11'b10101000100) ? 46'b0100111010011111011111001001110100111110111110 :
(key == 11'b10101000101) ? 46'b0100111001111111101111001001110011111111011110 :
(key == 11'b10101000110) ? 46'b0100111001100000000001101001110011000000000011 :
(key == 11'b10101000111) ? 46'b0100111001000000010111001001110010000000101110 :
(key == 11'b10101001000) ? 46'b0100111000100000101110001001110001000001011100 :
(key == 11'b10101001001) ? 46'b0100111000000001000110101001110000000010001101 :
(key == 11'b10101001010) ? 46'b0100110111100001100010001001101111000011000100 :
(key == 11'b10101001011) ? 46'b0100110111000010000000101001101110000100000001 :
(key == 11'b10101001100) ? 46'b0100110110100010100000101001101101000101000001 :
(key == 11'b10101001101) ? 46'b0100110110000011000010001001101100000110000100 :
(key == 11'b10101001110) ? 46'b0100110101100011100111101001101011000111001111 :
(key == 11'b10101001111) ? 46'b0100110101000100001110101001101010001000011101 :
(key == 11'b10101010000) ? 46'b0100110100100100110110101001101001001001101101 :
(key == 11'b10101010001) ? 46'b0100110100000101100010001001101000001011000100 :
(key == 11'b10101010010) ? 46'b0100110011100110001111101001100111001100011111 :
(key == 11'b10101010011) ? 46'b0100110011000110111111001001100110001101111110 :
(key == 11'b10101010100) ? 46'b0100110010100111110000101001100101001111100001 :
(key == 11'b10101010101) ? 46'b0100110010001000100100101001100100010001001001 :
(key == 11'b10101010110) ? 46'b0100110001101001011011001001100011010010110110 :
(key == 11'b10101010111) ? 46'b0100110001001010010011101001100010010100100111 :
(key == 11'b10101011000) ? 46'b0100110000101011001110001001100001010110011100 :
(key == 11'b10101011001) ? 46'b0100110000001100001010001001100000011000010100 :
(key == 11'b10101011010) ? 46'b0100101111101101001001101001011111011010010011 :
(key == 11'b10101011011) ? 46'b0100101111001110001010001001011110011100010100 :
(key == 11'b10101011100) ? 46'b0100101110101111001101101001011101011110011011 :
(key == 11'b10101011101) ? 46'b0100101110010000010011001001011100100000100110 :
(key == 11'b10101011110) ? 46'b0100101101110001011010001001011011100010110100 :
(key == 11'b10101011111) ? 46'b0100101101010010100100001001011010100101001000 :
(key == 11'b10101100000) ? 46'b0100101100110011110000001001011001100111100000 :
(key == 11'b10101100001) ? 46'b0100101100010100111101101001011000101001111011 :
(key == 11'b10101100010) ? 46'b0100101011110110001110001001010111101100011100 :
(key == 11'b10101100011) ? 46'b0100101011010111100000101001010110101111000001 :
(key == 11'b10101100100) ? 46'b0100101010111000110100101001010101110001101001 :
(key == 11'b10101100101) ? 46'b0100101010011010001011001001010100110100010110 :
(key == 11'b10101100110) ? 46'b0100101001111011100100001001010011110111001000 :
(key == 11'b10101100111) ? 46'b0100101001011100111111001001010010111001111110 :
(key == 11'b10101101000) ? 46'b0100101000111110011011001001010001111100110110 :
(key == 11'b10101101001) ? 46'b0100101000011111111010001001010000111111110100 :
(key == 11'b10101101010) ? 46'b0100101000000001011011001001010000000010110110 :
(key == 11'b10101101011) ? 46'b0100100111100010111111001001001111000101111110 :
(key == 11'b10101101100) ? 46'b0100100111000100100100001001001110001001001000 :
(key == 11'b10101101101) ? 46'b0100100110100110001100001001001101001100011000 :
(key == 11'b10101101110) ? 46'b0100100110000111110101001001001100001111101010 :
(key == 11'b10101101111) ? 46'b0100100101101001100001001001001011010011000010 :
(key == 11'b10101110000) ? 46'b0100100101001011001111001001001010010110011110 :
(key == 11'b10101110001) ? 46'b0100100100101100111110001001001001011001111100 :
(key == 11'b10101110010) ? 46'b0100100100001110110000101001001000011101100001 :
(key == 11'b10101110011) ? 46'b0100100011110000100100001001000111100001001000 :
(key == 11'b10101110100) ? 46'b0100100011010010011011001001000110100100110110 :
(key == 11'b10101110101) ? 46'b0100100010110100010010101001000101101000100101 :
(key == 11'b10101110110) ? 46'b0100100010010110001100001001000100101100011000 :
(key == 11'b10101110111) ? 46'b0100100001111000001001001001000011110000010010 :
(key == 11'b10101111000) ? 46'b0100100001011010000111001001000010110100001110 :
(key == 11'b10101111001) ? 46'b0100100000111100000111101001000001111000001111 :
(key == 11'b10101111010) ? 46'b0100100000011110001010001001000000111100010100 :
(key == 11'b10101111011) ? 46'b0100100000000000001110101001000000000000011101 :
(key == 11'b10101111100) ? 46'b0100011111100010010101001000111111000100101010 :
(key == 11'b10101111101) ? 46'b0100011111000100011110001000111110001000111100 :
(key == 11'b10101111110) ? 46'b0100011110100110101000101000111101001101010001 :
(key == 11'b10101111111) ? 46'b0100011110001000110101001000111100010001101010 :
(key == 11'b10110000000) ? 46'b0100011101101011000011001000111011010110000110 :
(key == 11'b10110000001) ? 46'b0100011101001101010100101000111010011010101001 :
(key == 11'b10110000010) ? 46'b0100011100101111100111001000111001011111001110 :
(key == 11'b10110000011) ? 46'b0100011100010001111100001000111000100011111000 :
(key == 11'b10110000100) ? 46'b0100011011110100010011001000110111101000100110 :
(key == 11'b10110000101) ? 46'b0100011011010110101011001000110110101101010110 :
(key == 11'b10110000110) ? 46'b0100011010111001000110001000110101110010001100 :
(key == 11'b10110000111) ? 46'b0100011010011011100011001000110100110111000110 :
(key == 11'b10110001000) ? 46'b0100011001111110000010001000110011111100000100 :
(key == 11'b10110001001) ? 46'b0100011001100000100011001000110011000001000110 :
(key == 11'b10110001010) ? 46'b0100011001000011000101101000110010000110001011 :
(key == 11'b10110001011) ? 46'b0100011000100101101010101000110001001011010101 :
(key == 11'b10110001100) ? 46'b0100011000001000010000101000110000010000100001 :
(key == 11'b10110001101) ? 46'b0100010111101010111001001000101111010101110010 :
(key == 11'b10110001110) ? 46'b0100010111001101100100001000101110011011001000 :
(key == 11'b10110001111) ? 46'b0100010110110000010001001000101101100000100010 :
(key == 11'b10110010000) ? 46'b0100010110010011000000001000101100100110000000 :
(key == 11'b10110010001) ? 46'b0100010101110101110000101000101011101011100001 :
(key == 11'b10110010010) ? 46'b0100010101011000100011101000101010110001000111 :
(key == 11'b10110010011) ? 46'b0100010100111011011000001000101001110110110000 :
(key == 11'b10110010100) ? 46'b0100010100011110001111001000101000111100011110 :
(key == 11'b10110010101) ? 46'b0100010100000001000111001000101000000010001110 :
(key == 11'b10110010110) ? 46'b0100010011100100000001001000100111001000000010 :
(key == 11'b10110010111) ? 46'b0100010011000110111110001000100110001101111100 :
(key == 11'b10110011000) ? 46'b0100010010101001111100101000100101010011111001 :
(key == 11'b10110011001) ? 46'b0100010010001100111100001000100100011001111000 :
(key == 11'b10110011010) ? 46'b0100010001101111111111001000100011011111111110 :
(key == 11'b10110011011) ? 46'b0100010001010011000011001000100010100110000110 :
(key == 11'b10110011100) ? 46'b0100010000110110001001001000100001101100010010 :
(key == 11'b10110011101) ? 46'b0100010000011001010001101000100000110010100011 :
(key == 11'b10110011110) ? 46'b0100001111111100011011001000011111111000110110 :
(key == 11'b10110011111) ? 46'b0100001111011111100111001000011110111111001110 :
(key == 11'b10110100000) ? 46'b0100001111000010110101001000011110000101101010 :
(key == 11'b10110100001) ? 46'b0100001110100110000101001000011101001100001010 :
(key == 11'b10110100010) ? 46'b0100001110001001010110001000011100010010101100 :
(key == 11'b10110100011) ? 46'b0100001101101100101010001000011011011001010100 :
(key == 11'b10110100100) ? 46'b0100001101001111111111101000011010011111111111 :
(key == 11'b10110100101) ? 46'b0100001100110011010111001000011001100110101110 :
(key == 11'b10110100110) ? 46'b0100001100010110110000101000011000101101100001 :
(key == 11'b10110100111) ? 46'b0100001011111010001011001000010111110100010110 :
(key == 11'b10110101000) ? 46'b0100001011011101101000101000010110111011010001 :
(key == 11'b10110101001) ? 46'b0100001011000001000111101000010110000010001111 :
(key == 11'b10110101010) ? 46'b0100001010100100101000101000010101001001010001 :
(key == 11'b10110101011) ? 46'b0100001010001000001011001000010100010000010110 :
(key == 11'b10110101100) ? 46'b0100001001101011110000001000010011010111100000 :
(key == 11'b10110101101) ? 46'b0100001001001111010110001000010010011110101100 :
(key == 11'b10110101110) ? 46'b0100001000110010111110101000010001100101111101 :
(key == 11'b10110101111) ? 46'b0100001000010110101001001000010000101101010010 :
(key == 11'b10110110000) ? 46'b0100000111111010010101001000001111110100101010 :
(key == 11'b10110110001) ? 46'b0100000111011110000011001000001110111100000110 :
(key == 11'b10110110010) ? 46'b0100000111000001110011001000001110000011100110 :
(key == 11'b10110110011) ? 46'b0100000110100101100100101000001101001011001001 :
(key == 11'b10110110100) ? 46'b0100000110001001011000001000001100010010110000 :
(key == 11'b10110110101) ? 46'b0100000101101101001101001000001011011010011010 :
(key == 11'b10110110110) ? 46'b0100000101010001000100101000001010100010001001 :
(key == 11'b10110110111) ? 46'b0100000100110100111101101000001001101001111011 :
(key == 11'b10110111000) ? 46'b0100000100011000111000101000001000110001110001 :
(key == 11'b10110111001) ? 46'b0100000011111100110110001000000111111001101100 :
(key == 11'b10110111010) ? 46'b0100000011100000110100001000000111000001101000 :
(key == 11'b10110111011) ? 46'b0100000011000100110101001000000110001001101010 :
(key == 11'b10110111100) ? 46'b0100000010101000110111101000000101010001101111 :
(key == 11'b10110111101) ? 46'b0100000010001100111011101000000100011001110111 :
(key == 11'b10110111110) ? 46'b0100000001110001000001001000000011100010000010 :
(key == 11'b10110111111) ? 46'b0100000001010101001001001000000010101010010010 :
(key == 11'b10111000000) ? 46'b0100000000111001010010001000000001110010100100 :
(key == 11'b10111000001) ? 46'b0100000000011101011110001000000000111010111100 :
(key == 11'b10111000010) ? 46'b0100000000000001101010101000000000000011010101 :
(key == 11'b10111000011) ? 46'b0011111111100101111010000111111111001011110100 :
(key == 11'b10111000100) ? 46'b0011111111001010001011000111111110010100010110 :
(key == 11'b10111000101) ? 46'b0011111110101110011101100111111101011100111011 :
(key == 11'b10111000110) ? 46'b0011111110010010110001100111111100100101100011 :
(key == 11'b10111000111) ? 46'b0011111101110111001000000111111011101110010000 :
(key == 11'b10111001000) ? 46'b0011111101011011100000100111111010110111000001 :
(key == 11'b10111001001) ? 46'b0011111100111111111010000111111001111111110100 :
(key == 11'b10111001010) ? 46'b0011111100100100010101100111111001001000101011 :
(key == 11'b10111001011) ? 46'b0011111100001000110010100111111000010001100101 :
(key == 11'b10111001100) ? 46'b0011111011101101010010000111110111011010100100 :
(key == 11'b10111001101) ? 46'b0011111011010001110011000111110110100011100110 :
(key == 11'b10111001110) ? 46'b0011111010110110010101100111110101101100101011 :
(key == 11'b10111001111) ? 46'b0011111010011010111010000111110100110101110100 :
(key == 11'b10111010000) ? 46'b0011111001111111100000000111110011111111000000 :
(key == 11'b10111010001) ? 46'b0011111001100100001000100111110011001000010001 :
(key == 11'b10111010010) ? 46'b0011111001001000110010000111110010010001100100 :
(key == 11'b10111010011) ? 46'b0011111000101101011101100111110001011010111011 :
(key == 11'b10111010100) ? 46'b0011111000010010001011000111110000100100010110 :
(key == 11'b10111010101) ? 46'b0011110111110110111010000111101111101101110100 :
(key == 11'b10111010110) ? 46'b0011110111011011101011000111101110110111010110 :
(key == 11'b10111010111) ? 46'b0011110111000000011101000111101110000000111010 :
(key == 11'b10111011000) ? 46'b0011110110100101010001000111101101001010100010 :
(key == 11'b10111011001) ? 46'b0011110110001010001000000111101100010100010000 :
(key == 11'b10111011010) ? 46'b0011110101101110111111100111101011011101111111 :
(key == 11'b10111011011) ? 46'b0011110101010011111001100111101010100111110011 :
(key == 11'b10111011100) ? 46'b0011110100111000110100000111101001110001101000 :
(key == 11'b10111011101) ? 46'b0011110100011101110001000111101000111011100010 :
(key == 11'b10111011110) ? 46'b0011110100000010110000100111101000000101100001 :
(key == 11'b10111011111) ? 46'b0011110011100111110000100111100111001111100001 :
(key == 11'b10111100000) ? 46'b0011110011001100110011000111100110011001100110 :
(key == 11'b10111100001) ? 46'b0011110010110001110110100111100101100011101101 :
(key == 11'b10111100010) ? 46'b0011110010010110111100000111100100101101111000 :
(key == 11'b10111100011) ? 46'b0011110001111100000011000111100011111000000110 :
(key == 11'b10111100100) ? 46'b0011110001100001001100100111100011000010011001 :
(key == 11'b10111100101) ? 46'b0011110001000110010111100111100010001100101111 :
(key == 11'b10111100110) ? 46'b0011110000101011100100000111100001010111001000 :
(key == 11'b10111100111) ? 46'b0011110000010000110010000111100000100001100100 :
(key == 11'b10111101000) ? 46'b0011101111110110000010000111011111101100000100 :
(key == 11'b10111101001) ? 46'b0011101111011011010011000111011110110110100110 :
(key == 11'b10111101010) ? 46'b0011101111000000100110000111011110000001001100 :
(key == 11'b10111101011) ? 46'b0011101110100101111011100111011101001011110111 :
(key == 11'b10111101100) ? 46'b0011101110001011010010000111011100010110100100 :
(key == 11'b10111101101) ? 46'b0011101101110000101011000111011011100001010110 :
(key == 11'b10111101110) ? 46'b0011101101010110000100100111011010101100001001 :
(key == 11'b10111101111) ? 46'b0011101100111011100000000111011001110111000000 :
(key == 11'b10111110000) ? 46'b0011101100100000111101000111011001000001111010 :
(key == 11'b10111110001) ? 46'b0011101100000110011100000111011000001100111000 :
(key == 11'b10111110010) ? 46'b0011101011101011111101000111010111010111111010 :
(key == 11'b10111110011) ? 46'b0011101011010001011111100111010110100010111111 :
(key == 11'b10111110100) ? 46'b0011101010110111000011000111010101101110000110 :
(key == 11'b10111110101) ? 46'b0011101010011100101001000111010100111001010010 :
(key == 11'b10111110110) ? 46'b0011101010000010010000000111010100000100100000 :
(key == 11'b10111110111) ? 46'b0011101001100111111010000111010011001111110100 :
(key == 11'b10111111000) ? 46'b0011101001001101100100000111010010011011001000 :
(key == 11'b10111111001) ? 46'b0011101000110011010000100111010001100110100001 :
(key == 11'b10111111010) ? 46'b0011101000011000111110000111010000110001111100 :
(key == 11'b10111111011) ? 46'b0011100111111110101110000111001111111101011100 :
(key == 11'b10111111100) ? 46'b0011100111100100011111100111001111001000111111 :
(key == 11'b10111111101) ? 46'b0011100111001010010010000111001110010100100100 :
(key == 11'b10111111110) ? 46'b0011100110110000000111000111001101100000001110 :
(key == 11'b10111111111) ? 46'b0011100110010101111101000111001100101011111010 :
(key == 11'b11000000000) ? 46'b0011100101111011110100100111001011110111101001 :
(key == 11'b11000000001) ? 46'b0011100101100001101110000111001011000011011100 :
(key == 11'b11000000010) ? 46'b0011100101000111101001100111001010001111010011 :
(key == 11'b11000000011) ? 46'b0011100100101101100110100111001001011011001101 :
(key == 11'b11000000100) ? 46'b0011100100010011100100000111001000100111001000 :
(key == 11'b11000000101) ? 46'b0011100011111001100011100111000111110011000111 :
(key == 11'b11000000110) ? 46'b0011100011011111100101100111000110111111001011 :
(key == 11'b11000000111) ? 46'b0011100011000101101001000111000110001011010010 :
(key == 11'b11000001000) ? 46'b0011100010101011101110000111000101010111011100 :
(key == 11'b11000001001) ? 46'b0011100010010001110100000111000100100011101000 :
(key == 11'b11000001010) ? 46'b0011100001110111111100000111000011101111111000 :
(key == 11'b11000001011) ? 46'b0011100001011110000110000111000010111100001100 :
(key == 11'b11000001100) ? 46'b0011100001000100010001000111000010001000100010 :
(key == 11'b11000001101) ? 46'b0011100000101010011101100111000001010100111011 :
(key == 11'b11000001110) ? 46'b0011100000010000101100100111000000100001011001 :
(key == 11'b11000001111) ? 46'b0011011111110110111100000110111111101101111000 :
(key == 11'b11000010000) ? 46'b0011011111011101001110000110111110111010011100 :
(key == 11'b11000010001) ? 46'b0011011111000011100001000110111110000111000010 :
(key == 11'b11000010010) ? 46'b0011011110101001110110000110111101010011101100 :
(key == 11'b11000010011) ? 46'b0011011110010000001100100110111100100000011001 :
(key == 11'b11000010100) ? 46'b0011011101110110100100100110111011101101001001 :
(key == 11'b11000010101) ? 46'b0011011101011100111101100110111010111001111011 :
(key == 11'b11000010110) ? 46'b0011011101000011011001000110111010000110110010 :
(key == 11'b11000010111) ? 46'b0011011100101001110101100110111001010011101011 :
(key == 11'b11000011000) ? 46'b0011011100010000010100000110111000100000101000 :
(key == 11'b11000011001) ? 46'b0011011011110110110011100110110111101101100111 :
(key == 11'b11000011010) ? 46'b0011011011011101010101000110110110111010101010 :
(key == 11'b11000011011) ? 46'b0011011011000011111000100110110110000111110001 :
(key == 11'b11000011100) ? 46'b0011011010101010011100100110110101010100111001 :
(key == 11'b11000011101) ? 46'b0011011010010001000010000110110100100010000100 :
(key == 11'b11000011110) ? 46'b0011011001110111101010100110110011101111010101 :
(key == 11'b11000011111) ? 46'b0011011001011110010011100110110010111100100111 :
(key == 11'b11000100000) ? 46'b0011011001000100111110000110110010001001111100 :
(key == 11'b11000100001) ? 46'b0011011000101011101010000110110001010111010100 :
(key == 11'b11000100010) ? 46'b0011011000010010011000000110110000100100110000 :
(key == 11'b11000100011) ? 46'b0011010111111001000111000110101111110010001110 :
(key == 11'b11000100100) ? 46'b0011010111011111111001000110101110111111110010 :
(key == 11'b11000100101) ? 46'b0011010111000110101011100110101110001101010111 :
(key == 11'b11000100110) ? 46'b0011010110101101011111100110101101011010111111 :
(key == 11'b11000100111) ? 46'b0011010110010100010100000110101100101000101000 :
(key == 11'b11000101000) ? 46'b0011010101111011001011100110101011110110010111 :
(key == 11'b11000101001) ? 46'b0011010101100010000100000110101011000100001000 :
(key == 11'b11000101010) ? 46'b0011010101001000111110000110101010010001111100 :
(key == 11'b11000101011) ? 46'b0011010100101111111001100110101001011111110011 :
(key == 11'b11000101100) ? 46'b0011010100010110110111000110101000101101101110 :
(key == 11'b11000101101) ? 46'b0011010011111101110110000110100111111011101100 :
(key == 11'b11000101110) ? 46'b0011010011100100110110000110100111001001101100 :
(key == 11'b11000101111) ? 46'b0011010011001011111000000110100110010111110000 :
(key == 11'b11000110000) ? 46'b0011010010110010111011000110100101100101110110 :
(key == 11'b11000110001) ? 46'b0011010010011010000000000110100100110100000000 :
(key == 11'b11000110010) ? 46'b0011010010000001000110000110100100000010001100 :
(key == 11'b11000110011) ? 46'b0011010001101000001101100110100011010000011011 :
(key == 11'b11000110100) ? 46'b0011010001001111010111000110100010011110101110 :
(key == 11'b11000110101) ? 46'b0011010000110110100001100110100001101101000011 :
(key == 11'b11000110110) ? 46'b0011010000011101101110000110100000111011011100 :
(key == 11'b11000110111) ? 46'b0011010000000100111011100110100000001001110111 :
(key == 11'b11000111000) ? 46'b0011001111101100001011000110011111011000010110 :
(key == 11'b11000111001) ? 46'b0011001111010011011100000110011110100110111000 :
(key == 11'b11000111010) ? 46'b0011001110111010101110100110011101110101011101 :
(key == 11'b11000111011) ? 46'b0011001110100010000010100110011101000100000101 :
(key == 11'b11000111100) ? 46'b0011001110001001010111000110011100010010101110 :
(key == 11'b11000111101) ? 46'b0011001101110000101101100110011011100001011011 :
(key == 11'b11000111110) ? 46'b0011001101011000000110000110011010110000001100 :
(key == 11'b11000111111) ? 46'b0011001100111111011111100110011001111110111111 :
(key == 11'b11001000000) ? 46'b0011001100100110111010100110011001001101110101 :
(key == 11'b11001000001) ? 46'b0011001100001110010111100110011000011100101111 :
(key == 11'b11001000010) ? 46'b0011001011110101110101100110010111101011101011 :
(key == 11'b11001000011) ? 46'b0011001011011101010101000110010110111010101010 :
(key == 11'b11001000100) ? 46'b0011001011000100110110000110010110001001101100 :
(key == 11'b11001000101) ? 46'b0011001010101100011000000110010101011000110000 :
(key == 11'b11001000110) ? 46'b0011001010010011111101000110010100100111111010 :
(key == 11'b11001000111) ? 46'b0011001001111011100010000110010011110111000100 :
(key == 11'b11001001000) ? 46'b0011001001100011001000100110010011000110010001 :
(key == 11'b11001001001) ? 46'b0011001001001010110001000110010010010101100010 :
(key == 11'b11001001010) ? 46'b0011001000110010011011000110010001100100110110 :
(key == 11'b11001001011) ? 46'b0011001000011010000110000110010000110100001100 :
(key == 11'b11001001100) ? 46'b0011001000000001110011000110010000000011100110 :
(key == 11'b11001001101) ? 46'b0011000111101001100001000110001111010011000010 :
(key == 11'b11001001110) ? 46'b0011000111010001010000100110001110100010100001 :
(key == 11'b11001001111) ? 46'b0011000110111001000001000110001101110010000010 :
(key == 11'b11001010000) ? 46'b0011000110100000110100000110001101000001101000 :
(key == 11'b11001010001) ? 46'b0011000110001000101000000110001100010001010000 :
(key == 11'b11001010010) ? 46'b0011000101110000011101000110001011100000111010 :
(key == 11'b11001010011) ? 46'b0011000101011000010100000110001010110000101000 :
(key == 11'b11001010100) ? 46'b0011000101000000001100000110001010000000011000 :
(key == 11'b11001010101) ? 46'b0011000100101000000110000110001001010000001100 :
(key == 11'b11001010110) ? 46'b0011000100010000000001000110001000100000000010 :
(key == 11'b11001010111) ? 46'b0011000011110111111100100110000111101111111001 :
(key == 11'b11001011000) ? 46'b0011000011011111111011000110000110111111110110 :
(key == 11'b11001011001) ? 46'b0011000011000111111010000110000110001111110100 :
(key == 11'b11001011010) ? 46'b0011000010101111111011000110000101011111110110 :
(key == 11'b11001011011) ? 46'b0011000010010111111101100110000100101111111011 :
(key == 11'b11001011100) ? 46'b0011000010000000000001000110000100000000000010 :
(key == 11'b11001011101) ? 46'b0011000001101000000101100110000011010000001011 :
(key == 11'b11001011110) ? 46'b0011000001010000001011100110000010100000010111 :
(key == 11'b11001011111) ? 46'b0011000000111000010100000110000001110000101000 :
(key == 11'b11001100000) ? 46'b0011000000100000011101000110000001000000111010 :
(key == 11'b11001100001) ? 46'b0011000000001000101000000110000000010001010000 :
(key == 11'b11001100010) ? 46'b0010111111110000110011100101111111100001100111 :
(key == 11'b11001100011) ? 46'b0010111111011001000000100101111110110010000001 :
(key == 11'b11001100100) ? 46'b0010111111000001001111100101111110000010011111 :
(key == 11'b11001100101) ? 46'b0010111110101001011111100101111101010010111111 :
(key == 11'b11001100110) ? 46'b0010111110010001110001000101111100100011100010 :
(key == 11'b11001100111) ? 46'b0010111101111010000100000101111011110100001000 :
(key == 11'b11001101000) ? 46'b0010111101100010011000000101111011000100110000 :
(key == 11'b11001101001) ? 46'b0010111101001010101110000101111010010101011100 :
(key == 11'b11001101010) ? 46'b0010111100110011000101000101111001100110001010 :
(key == 11'b11001101011) ? 46'b0010111100011011011101100101111000110110111011 :
(key == 11'b11001101100) ? 46'b0010111100000011111000000101111000000111110000 :
(key == 11'b11001101101) ? 46'b0010111011101100010011000101110111011000100110 :
(key == 11'b11001101110) ? 46'b0010111011010100110000000101110110101001100000 :
(key == 11'b11001101111) ? 46'b0010111010111101001110000101110101111010011100 :
(key == 11'b11001110000) ? 46'b0010111010100101101100100101110101001011011001 :
(key == 11'b11001110001) ? 46'b0010111010001110001101100101110100011100011011 :
(key == 11'b11001110010) ? 46'b0010111001110110101111100101110011101101011111 :
(key == 11'b11001110011) ? 46'b0010111001011111010011000101110010111110100110 :
(key == 11'b11001110100) ? 46'b0010111001000111111000100101110010001111110001 :
(key == 11'b11001110101) ? 46'b0010111000110000011110000101110001100000111100 :
(key == 11'b11001110110) ? 46'b0010111000011001000101000101110000110010001010 :
(key == 11'b11001110111) ? 46'b0010111000000001101110100101110000000011011101 :
(key == 11'b11001111000) ? 46'b0010110111101010011001000101101111010100110010 :
(key == 11'b11001111001) ? 46'b0010110111010011000101000101101110100110001010 :
(key == 11'b11001111010) ? 46'b0010110110111011110001100101101101110111100011 :
(key == 11'b11001111011) ? 46'b0010110110100100011111000101101101001000111110 :
(key == 11'b11001111100) ? 46'b0010110110001101001111000101101100011010011110 :
(key == 11'b11001111101) ? 46'b0010110101110110000000000101101011101100000000 :
(key == 11'b11001111110) ? 46'b0010110101011110110010100101101010111101100101 :
(key == 11'b11001111111) ? 46'b0010110101000111100110000101101010001111001100 :
(key == 11'b11010000000) ? 46'b0010110100110000011011100101101001100000110111 :
(key == 11'b11010000001) ? 46'b0010110100011001010001100101101000110010100011 :
(key == 11'b11010000010) ? 46'b0010110100000010001001000101101000000100010010 :
(key == 11'b11010000011) ? 46'b0010110011101011000010000101100111010110000100 :
(key == 11'b11010000100) ? 46'b0010110011010011111100000101100110100111111000 :
(key == 11'b11010000101) ? 46'b0010110010111100111000000101100101111001110000 :
(key == 11'b11010000110) ? 46'b0010110010100101110101000101100101001011101010 :
(key == 11'b11010000111) ? 46'b0010110010001110110100000101100100011101101000 :
(key == 11'b11010001000) ? 46'b0010110001110111110011000101100011101111100110 :
(key == 11'b11010001001) ? 46'b0010110001100000110100000101100011000001101000 :
(key == 11'b11010001010) ? 46'b0010110001001001110110100101100010010011101101 :
(key == 11'b11010001011) ? 46'b0010110000110010111010000101100001100101110100 :
(key == 11'b11010001100) ? 46'b0010110000011011111110100101100000110111111101 :
(key == 11'b11010001101) ? 46'b0010110000000101000101000101100000001010001010 :
(key == 11'b11010001110) ? 46'b0010101111101110001100100101011111011100011001 :
(key == 11'b11010001111) ? 46'b0010101111010111010101000101011110101110101010 :
(key == 11'b11010010000) ? 46'b0010101111000000100000000101011110000001000000 :
(key == 11'b11010010001) ? 46'b0010101110101001101011000101011101010011010110 :
(key == 11'b11010010010) ? 46'b0010101110010010110111100101011100100101101111 :
(key == 11'b11010010011) ? 46'b0010101101111100000101100101011011111000001011 :
(key == 11'b11010010100) ? 46'b0010101101100101010101000101011011001010101010 :
(key == 11'b11010010101) ? 46'b0010101101001110100110000101011010011101001100 :
(key == 11'b11010010110) ? 46'b0010101100110111110111100101011001101111101111 :
(key == 11'b11010010111) ? 46'b0010101100100001001011000101011001000010010110 :
(key == 11'b11010011000) ? 46'b0010101100001010011111100101011000010100111111 :
(key == 11'b11010011001) ? 46'b0010101011110011110101000101010111100111101010 :
(key == 11'b11010011010) ? 46'b0010101011011101001100000101010110111010011000 :
(key == 11'b11010011011) ? 46'b0010101011000110100101000101010110001101001010 :
(key == 11'b11010011100) ? 46'b0010101010101111111110000101010101011111111100 :
(key == 11'b11010011101) ? 46'b0010101010011001011001100101010100110010110011 :
(key == 11'b11010011110) ? 46'b0010101010000010110101100101010100000101101011 :
(key == 11'b11010011111) ? 46'b0010101001101100010010100101010011011000100101 :
(key == 11'b11010100000) ? 46'b0010101001010101110001100101010010101011100011 :
(key == 11'b11010100001) ? 46'b0010101000111111010010000101010001111110100100 :
(key == 11'b11010100010) ? 46'b0010101000101000110011000101010001010001100110 :
(key == 11'b11010100011) ? 46'b0010101000010010010101000101010000100100101010 :
(key == 11'b11010100100) ? 46'b0010100111111011111001000101001111110111110010 :
(key == 11'b11010100101) ? 46'b0010100111100101011110100101001111001010111101 :
(key == 11'b11010100110) ? 46'b0010100111001111000101000101001110011110001010 :
(key == 11'b11010100111) ? 46'b0010100110111000101100100101001101110001011001 :
(key == 11'b11010101000) ? 46'b0010100110100010010101100101001101000100101011 :
(key == 11'b11010101001) ? 46'b0010100110001011111111100101001100010111111111 :
(key == 11'b11010101010) ? 46'b0010100101110101101011000101001011101011010110 :
(key == 11'b11010101011) ? 46'b0010100101011111011000000101001010111110110000 :
(key == 11'b11010101100) ? 46'b0010100101001001000101100101001010010010001011 :
(key == 11'b11010101101) ? 46'b0010100100110010110101000101001001100101101010 :
(key == 11'b11010101110) ? 46'b0010100100011100100101100101001000111001001011 :
(key == 11'b11010101111) ? 46'b0010100100000110010111000101001000001100101110 :
(key == 11'b11010110000) ? 46'b0010100011110000001010000101000111100000010100 :
(key == 11'b11010110001) ? 46'b0010100011011001111110000101000110110011111100 :
(key == 11'b11010110010) ? 46'b0010100011000011110011100101000110000111100111 :
(key == 11'b11010110011) ? 46'b0010100010101101101010000101000101011011010100 :
(key == 11'b11010110100) ? 46'b0010100010010111100010000101000100101111000100 :
(key == 11'b11010110101) ? 46'b0010100010000001011011000101000100000010110110 :
(key == 11'b11010110110) ? 46'b0010100001101011010101100101000011010110101011 :
(key == 11'b11010110111) ? 46'b0010100001010101010001000101000010101010100010 :
(key == 11'b11010111000) ? 46'b0010100000111111001110000101000001111110011100 :
(key == 11'b11010111001) ? 46'b0010100000101001001100000101000001010010011000 :
(key == 11'b11010111010) ? 46'b0010100000010011001011000101000000100110010110 :
(key == 11'b11010111011) ? 46'b0010011111111101001100000100111111111010011000 :
(key == 11'b11010111100) ? 46'b0010011111100111001101000100111111001110011010 :
(key == 11'b11010111101) ? 46'b0010011111010001010000100100111110100010100001 :
(key == 11'b11010111110) ? 46'b0010011110111011010100100100111101110110101001 :
(key == 11'b11010111111) ? 46'b0010011110100101011010100100111101001010110101 :
(key == 11'b11011000000) ? 46'b0010011110001111100001100100111100011111000011 :
(key == 11'b11011000001) ? 46'b0010011101111001101001000100111011110011010010 :
(key == 11'b11011000010) ? 46'b0010011101100011110001000100111011000111100010 :
(key == 11'b11011000011) ? 46'b0010011101001101111011100100111010011011110111 :
(key == 11'b11011000100) ? 46'b0010011100111000000111100100111001110000001111 :
(key == 11'b11011000101) ? 46'b0010011100100010010100000100111001000100101000 :
(key == 11'b11011000110) ? 46'b0010011100001100100010000100111000011001000100 :
(key == 11'b11011000111) ? 46'b0010011011110110110001000100110111101101100010 :
(key == 11'b11011001000) ? 46'b0010011011100001000001100100110111000010000011 :
(key == 11'b11011001001) ? 46'b0010011011001011010011000100110110010110100110 :
(key == 11'b11011001010) ? 46'b0010011010110101100101100100110101101011001011 :
(key == 11'b11011001011) ? 46'b0010011010011111111001100100110100111111110011 :
(key == 11'b11011001100) ? 46'b0010011010001010001110000100110100010100011100 :
(key == 11'b11011001101) ? 46'b0010011001110100100100100100110011101001001001 :
(key == 11'b11011001110) ? 46'b0010011001011110111100100100110010111101111001 :
(key == 11'b11011001111) ? 46'b0010011001001001010101100100110010010010101011 :
(key == 11'b11011010000) ? 46'b0010011000110011101111000100110001100111011110 :
(key == 11'b11011010001) ? 46'b0010011000011110001010100100110000111100010101 :
(key == 11'b11011010010) ? 46'b0010011000001000100110100100110000010001001101 :
(key == 11'b11011010011) ? 46'b0010010111110011000011100100101111100110000111 :
(key == 11'b11011010100) ? 46'b0010010111011101100010000100101110111011000100 :
(key == 11'b11011010101) ? 46'b0010010111001000000010000100101110010000000100 :
(key == 11'b11011010110) ? 46'b0010010110110010100011000100101101100101000110 :
(key == 11'b11011010111) ? 46'b0010010110011101000101000100101100111010001010 :
(key == 11'b11011011000) ? 46'b0010010110000111101000100100101100001111010001 :
(key == 11'b11011011001) ? 46'b0010010101110010001101000100101011100100011010 :
(key == 11'b11011011010) ? 46'b0010010101011100110011000100101010111001100110 :
(key == 11'b11011011011) ? 46'b0010010101000111011001000100101010001110110010 :
(key == 11'b11011011100) ? 46'b0010010100110010000001000100101001100100000010 :
(key == 11'b11011011101) ? 46'b0010010100011100101010100100101000111001010101 :
(key == 11'b11011011110) ? 46'b0010010100000111010100100100101000001110101001 :
(key == 11'b11011011111) ? 46'b0010010011110010000001000100100111100100000010 :
(key == 11'b11011100000) ? 46'b0010010011011100101101000100100110111001011010 :
(key == 11'b11011100001) ? 46'b0010010011000111011011000100100110001110110110 :
(key == 11'b11011100010) ? 46'b0010010010110010001010000100100101100100010100 :
(key == 11'b11011100011) ? 46'b0010010010011100111010000100100100111001110100 :
(key == 11'b11011100100) ? 46'b0010010010000111101011100100100100001111010111 :
(key == 11'b11011100101) ? 46'b0010010001110010011110000100100011100100111100 :
(key == 11'b11011100110) ? 46'b0010010001011101010001100100100010111010100011 :
(key == 11'b11011100111) ? 46'b0010010001001000000110000100100010010000001100 :
(key == 11'b11011101000) ? 46'b0010010000110010111100000100100001100101111000 :
(key == 11'b11011101001) ? 46'b0010010000011101110011000100100000111011100110 :
(key == 11'b11011101010) ? 46'b0010010000001000101011000100100000010001010110 :
(key == 11'b11011101011) ? 46'b0010001111110011100100100100011111100111001001 :
(key == 11'b11011101100) ? 46'b0010001111011110011111000100011110111100111110 :
(key == 11'b11011101101) ? 46'b0010001111001001011011000100011110010010110110 :
(key == 11'b11011101110) ? 46'b0010001110110100010111100100011101101000101111 :
(key == 11'b11011101111) ? 46'b0010001110011111010101000100011100111110101010 :
(key == 11'b11011110000) ? 46'b0010001110001010010100000100011100010100101000 :
(key == 11'b11011110001) ? 46'b0010001101110101010100000100011011101010101000 :
(key == 11'b11011110010) ? 46'b0010001101100000010110000100011011000000101100 :
(key == 11'b11011110011) ? 46'b0010001101001011011001000100011010010110110010 :
(key == 11'b11011110100) ? 46'b0010001100110110011100000100011001101100111000 :
(key == 11'b11011110101) ? 46'b0010001100100001100000100100011001000011000001 :
(key == 11'b11011110110) ? 46'b0010001100001100100110100100011000011001001101 :
(key == 11'b11011110111) ? 46'b0010001011110111101110000100010111101111011100 :
(key == 11'b11011111000) ? 46'b0010001011100010110101100100010111000101101011 :
(key == 11'b11011111001) ? 46'b0010001011001101111111000100010110011011111110 :
(key == 11'b11011111010) ? 46'b0010001010111001001001000100010101110010010010 :
(key == 11'b11011111011) ? 46'b0010001010100100010100100100010101001000101001 :
(key == 11'b11011111100) ? 46'b0010001010001111100001000100010100011111000010 :
(key == 11'b11011111101) ? 46'b0010001001111010101111000100010011110101011110 :
(key == 11'b11011111110) ? 46'b0010001001100101111101100100010011001011111011 :
(key == 11'b11011111111) ? 46'b0010001001010001001101000100010010100010011010 :
(key == 11'b11100000000) ? 46'b0010001000111100011110000100010001111000111100 :
(key == 11'b11100000001) ? 46'b0010001000100111110000000100010001001111100000 :
(key == 11'b11100000010) ? 46'b0010001000010011000100000100010000100110001000 :
(key == 11'b11100000011) ? 46'b0010000111111110011000000100001111111100110000 :
(key == 11'b11100000100) ? 46'b0010000111101001101110000100001111010011011100 :
(key == 11'b11100000101) ? 46'b0010000111010101000100100100001110101010001001 :
(key == 11'b11100000110) ? 46'b0010000111000000011100000100001110000000111000 :
(key == 11'b11100000111) ? 46'b0010000110101011110100100100001101010111101001 :
(key == 11'b11100001000) ? 46'b0010000110010111001110100100001100101110011101 :
(key == 11'b11100001001) ? 46'b0010000110000010101001000100001100000101010010 :
(key == 11'b11100001010) ? 46'b0010000101101110000101000100001011011100001010 :
(key == 11'b11100001011) ? 46'b0010000101011001100010100100001010110011000101 :
(key == 11'b11100001100) ? 46'b0010000101000101000001000100001010001010000010 :
(key == 11'b11100001101) ? 46'b0010000100110000100000100100001001100001000001 :
(key == 11'b11100001110) ? 46'b0010000100011100000000000100001000111000000000 :
(key == 11'b11100001111) ? 46'b0010000100000111100010000100001000001111000100 :
(key == 11'b11100010000) ? 46'b0010000011110011000100100100000111100110001001 :
(key == 11'b11100010001) ? 46'b0010000011011110101001000100000110111101010010 :
(key == 11'b11100010010) ? 46'b0010000011001010001101000100000110010100011010 :
(key == 11'b11100010011) ? 46'b0010000010110101110011000100000101101011100110 :
(key == 11'b11100010100) ? 46'b0010000010100001011010000100000101000010110100 :
(key == 11'b11100010101) ? 46'b0010000010001101000010000100000100011010000100 :
(key == 11'b11100010110) ? 46'b0010000001111000101011000100000011110001010110 :
(key == 11'b11100010111) ? 46'b0010000001100100010101000100000011001000101010 :
(key == 11'b11100011000) ? 46'b0010000001010000000000100100000010100000000001 :
(key == 11'b11100011001) ? 46'b0010000000111011101101000100000001110111011010 :
(key == 11'b11100011010) ? 46'b0010000000100111011010000100000001001110110100 :
(key == 11'b11100011011) ? 46'b0010000000010011001001000100000000100110010010 :
(key == 11'b11100011100) ? 46'b0001111111111110111000100011111111111101110001 :
(key == 11'b11100011101) ? 46'b0001111111101010101001000011111111010101010010 :
(key == 11'b11100011110) ? 46'b0001111111010110011010100011111110101100110101 :
(key == 11'b11100011111) ? 46'b0001111111000010001101000011111110000100011010 :
(key == 11'b11100100000) ? 46'b0001111110101110000000100011111101011100000001 :
(key == 11'b11100100001) ? 46'b0001111110011001110110000011111100110011101100 :
(key == 11'b11100100010) ? 46'b0001111110000101101011100011111100001011010111 :
(key == 11'b11100100011) ? 46'b0001111101110001100010000011111011100011000100 :
(key == 11'b11100100100) ? 46'b0001111101011101011011000011111010111010110110 :
(key == 11'b11100100101) ? 46'b0001111101001001010100000011111010010010101000 :
(key == 11'b11100100110) ? 46'b0001111100110101001110000011111001101010011100 :
(key == 11'b11100100111) ? 46'b0001111100100001001001000011111001000010010010 :
(key == 11'b11100101000) ? 46'b0001111100001101000101100011111000011010001011 :
(key == 11'b11100101001) ? 46'b0001111011111001000011000011110111110010000110 :
(key == 11'b11100101010) ? 46'b0001111011100101000001000011110111001010000010 :
(key == 11'b11100101011) ? 46'b0001111011010001000000100011110110100010000001 :
(key == 11'b11100101100) ? 46'b0001111010111101000000100011110101111010000001 :
(key == 11'b11100101101) ? 46'b0001111010101001000010100011110101010010000101 :
(key == 11'b11100101110) ? 46'b0001111010010101000101000011110100101010001010 :
(key == 11'b11100101111) ? 46'b0001111010000001001000100011110100000010010001 :
(key == 11'b11100110000) ? 46'b0001111001101101001101000011110011011010011010 :
(key == 11'b11100110001) ? 46'b0001111001011001010011000011110010110010100110 :
(key == 11'b11100110010) ? 46'b0001111001000101011001000011110010001010110010 :
(key == 11'b11100110011) ? 46'b0001111000110001100001000011110001100011000010 :
(key == 11'b11100110100) ? 46'b0001111000011101101010000011110000111011010100 :
(key == 11'b11100110101) ? 46'b0001111000001001110100000011110000010011101000 :
(key == 11'b11100110110) ? 46'b0001110111110101111110000011101111101011111100 :
(key == 11'b11100110111) ? 46'b0001110111100010001010000011101111000100010100 :
(key == 11'b11100111000) ? 46'b0001110111001110010111000011101110011100101110 :
(key == 11'b11100111001) ? 46'b0001110110111010100101000011101101110101001010 :
(key == 11'b11100111010) ? 46'b0001110110100110110100000011101101001101101000 :
(key == 11'b11100111011) ? 46'b0001110110010011000100000011101100100110001000 :
(key == 11'b11100111100) ? 46'b0001110101111111010101000011101011111110101010 :
(key == 11'b11100111101) ? 46'b0001110101101011100110100011101011010111001101 :
(key == 11'b11100111110) ? 46'b0001110101010111111001100011101010101111110011 :
(key == 11'b11100111111) ? 46'b0001110101000100001101100011101010001000011011 :
(key == 11'b11101000000) ? 46'b0001110100110000100011000011101001100001000110 :
(key == 11'b11101000001) ? 46'b0001110100011100111001100011101000111001110011 :
(key == 11'b11101000010) ? 46'b0001110100001001010000000011101000010010100000 :
(key == 11'b11101000011) ? 46'b0001110011110101101000000011100111101011010000 :
(key == 11'b11101000100) ? 46'b0001110011100010000001000011100111000100000010 :
(key == 11'b11101000101) ? 46'b0001110011001110011011100011100110011100110111 :
(key == 11'b11101000110) ? 46'b0001110010111010110110100011100101110101101101 :
(key == 11'b11101000111) ? 46'b0001110010100111010011000011100101001110100110 :
(key == 11'b11101001000) ? 46'b0001110010010011110000000011100100100111100000 :
(key == 11'b11101001001) ? 46'b0001110010000000001110000011100100000000011100 :
(key == 11'b11101001010) ? 46'b0001110001101100101101100011100011011001011011 :
(key == 11'b11101001011) ? 46'b0001110001011001001101000011100010110010011010 :
(key == 11'b11101001100) ? 46'b0001110001000101101111000011100010001011011110 :
(key == 11'b11101001101) ? 46'b0001110000110010010000100011100001100100100001 :
(key == 11'b11101001110) ? 46'b0001110000011110110100000011100000111101101000 :
(key == 11'b11101001111) ? 46'b0001110000001011011000100011100000010110110001 :
(key == 11'b11101010000) ? 46'b0001101111110111111101100011011111101111111011 :
(key == 11'b11101010001) ? 46'b0001101111100100100011100011011111001001000111 :
(key == 11'b11101010010) ? 46'b0001101111010001001010100011011110100010010101 :
(key == 11'b11101010011) ? 46'b0001101110111101110010100011011101111011100101 :
(key == 11'b11101010100) ? 46'b0001101110101010011100000011011101010100111000 :
(key == 11'b11101010101) ? 46'b0001101110010111000110000011011100101110001100 :
(key == 11'b11101010110) ? 46'b0001101110000011110001000011011100000111100010 :
(key == 11'b11101010111) ? 46'b0001101101110000011101100011011011100000111011 :
(key == 11'b11101011000) ? 46'b0001101101011101001010100011011010111010010101 :
(key == 11'b11101011001) ? 46'b0001101101001001111001000011011010010011110010 :
(key == 11'b11101011010) ? 46'b0001101100110110101000000011011001101101010000 :
(key == 11'b11101011011) ? 46'b0001101100100011010111100011011001000110101111 :
(key == 11'b11101011100) ? 46'b0001101100010000001001000011011000100000010010 :
(key == 11'b11101011101) ? 46'b0001101011111100111010100011010111111001110101 :
(key == 11'b11101011110) ? 46'b0001101011101001101101000011010111010011011010 :
(key == 11'b11101011111) ? 46'b0001101011010110100001100011010110101101000011 :
(key == 11'b11101100000) ? 46'b0001101011000011010111000011010110000110101110 :
(key == 11'b11101100001) ? 46'b0001101010110000001100100011010101100000011001 :
(key == 11'b11101100010) ? 46'b0001101010011101000011100011010100111010000111 :
(key == 11'b11101100011) ? 46'b0001101010001001111011100011010100010011110111 :
(key == 11'b11101100100) ? 46'b0001101001110110110100000011010011101101101000 :
(key == 11'b11101100101) ? 46'b0001101001100011101110000011010011000111011100 :
(key == 11'b11101100110) ? 46'b0001101001010000101000100011010010100001010001 :
(key == 11'b11101100111) ? 46'b0001101000111101100100000011010001111011001000 :
(key == 11'b11101101000) ? 46'b0001101000101010100001000011010001010101000010 :
(key == 11'b11101101001) ? 46'b0001101000010111011110100011010000101110111101 :
(key == 11'b11101101010) ? 46'b0001101000000100011101000011010000001000111010 :
(key == 11'b11101101011) ? 46'b0001100111110001011100100011001111100010111001 :
(key == 11'b11101101100) ? 46'b0001100111011110011101000011001110111100111010 :
(key == 11'b11101101101) ? 46'b0001100111001011011110100011001110010110111101 :
(key == 11'b11101101110) ? 46'b0001100110111000100001000011001101110001000010 :
(key == 11'b11101101111) ? 46'b0001100110100101100100100011001101001011001001 :
(key == 11'b11101110000) ? 46'b0001100110010010101001000011001100100101010010 :
(key == 11'b11101110001) ? 46'b0001100101111111101110000011001011111111011100 :
(key == 11'b11101110010) ? 46'b0001100101101100110101000011001011011001101010 :
(key == 11'b11101110011) ? 46'b0001100101011001111100000011001010110011111000 :
(key == 11'b11101110100) ? 46'b0001100101000111000100000011001010001110001000 :
(key == 11'b11101110101) ? 46'b0001100100110100001101000011001001101000011010 :
(key == 11'b11101110110) ? 46'b0001100100100001010111000011001001000010101110 :
(key == 11'b11101110111) ? 46'b0001100100001110100010000011001000011101000100 :
(key == 11'b11101111000) ? 46'b0001100011111011101110000011000111110111011100 :
(key == 11'b11101111001) ? 46'b0001100011101000111011000011000111010001110110 :
(key == 11'b11101111010) ? 46'b0001100011010110001001000011000110101100010010 :
(key == 11'b11101111011) ? 46'b0001100011000011011000000011000110000110110000 :
(key == 11'b11101111100) ? 46'b0001100010110000100111000011000101100001001110 :
(key == 11'b11101111101) ? 46'b0001100010011101111000000011000100111011110000 :
(key == 11'b11101111110) ? 46'b0001100010001011001010000011000100010110010100 :
(key == 11'b11101111111) ? 46'b0001100001111000011100100011000011110000111001 :
(key == 11'b11110000000) ? 46'b0001100001100101110000000011000011001011100000 :
(key == 11'b11110000001) ? 46'b0001100001010011000100000011000010100110001000 :
(key == 11'b11110000010) ? 46'b0001100001000000011001100011000010000000110011 :
(key == 11'b11110000011) ? 46'b0001100000101101110000000011000001011011100000 :
(key == 11'b11110000100) ? 46'b0001100000011011000111000011000000110110001110 :
(key == 11'b11110000101) ? 46'b0001100000001000011111000011000000010000111110 :
(key == 11'b11110000110) ? 46'b0001011111110101111001000010111111101011110010 :
(key == 11'b11110000111) ? 46'b0001011111100011010010100010111111000110100101 :
(key == 11'b11110001000) ? 46'b0001011111010000101101100010111110100001011011 :
(key == 11'b11110001001) ? 46'b0001011110111110001001000010111101111100010010 :
(key == 11'b11110001010) ? 46'b0001011110101011100110000010111101010111001100 :
(key == 11'b11110001011) ? 46'b0001011110011001000011100010111100110010000111 :
(key == 11'b11110001100) ? 46'b0001011110000110100010000010111100001101000100 :
(key == 11'b11110001101) ? 46'b0001011101110100000001100010111011101000000011 :
(key == 11'b11110001110) ? 46'b0001011101100001100010000010111011000011000100 :
(key == 11'b11110001111) ? 46'b0001011101001111000011100010111010011110000111 :
(key == 11'b11110010000) ? 46'b0001011100111100100110000010111001111001001100 :
(key == 11'b11110010001) ? 46'b0001011100101010001001000010111001010100010010 :
(key == 11'b11110010010) ? 46'b0001011100010111101101000010111000101111011010 :
(key == 11'b11110010011) ? 46'b0001011100000101010010000010111000001010100100 :
(key == 11'b11110010100) ? 46'b0001011011110010110111100010110111100101101111 :
(key == 11'b11110010101) ? 46'b0001011011100000011111000010110111000000111110 :
(key == 11'b11110010110) ? 46'b0001011011001110000111000010110110011100001110 :
(key == 11'b11110010111) ? 46'b0001011010111011101111000010110101110111011110 :
(key == 11'b11110011000) ? 46'b0001011010101001011001000010110101010010110010 :
(key == 11'b11110011001) ? 46'b0001011010010111000100000010110100101110001000 :
(key == 11'b11110011010) ? 46'b0001011010000100101110100010110100001001011101 :
(key == 11'b11110011011) ? 46'b0001011001110010011011000010110011100100110110 :
(key == 11'b11110011100) ? 46'b0001011001100000001000100010110011000000010001 :
(key == 11'b11110011101) ? 46'b0001011001001101110110100010110010011011101101 :
(key == 11'b11110011110) ? 46'b0001011000111011100101000010110001110111001010 :
(key == 11'b11110011111) ? 46'b0001011000101001010101000010110001010010101010 :
(key == 11'b11110100000) ? 46'b0001011000010111000110000010110000101110001100 :
(key == 11'b11110100001) ? 46'b0001011000000100110111100010110000001001101111 :
(key == 11'b11110100010) ? 46'b0001010111110010101010100010101111100101010101 :
(key == 11'b11110100011) ? 46'b0001010111100000011101100010101111000000111011 :
(key == 11'b11110100100) ? 46'b0001010111001110010001100010101110011100100011 :
(key == 11'b11110100101) ? 46'b0001010110111100000111000010101101111000001110 :
(key == 11'b11110100110) ? 46'b0001010110101001111110000010101101010011111100 :
(key == 11'b11110100111) ? 46'b0001010110010111110100100010101100101111101001 :
(key == 11'b11110101000) ? 46'b0001010110000101101100000010101100001011011000 :
(key == 11'b11110101001) ? 46'b0001010101110011100101100010101011100111001011 :
(key == 11'b11110101010) ? 46'b0001010101100001011111000010101011000010111110 :
(key == 11'b11110101011) ? 46'b0001010101001111011001100010101010011110110011 :
(key == 11'b11110101100) ? 46'b0001010100111101010101000010101001111010101010 :
(key == 11'b11110101101) ? 46'b0001010100101011010001000010101001010110100010 :
(key == 11'b11110101110) ? 46'b0001010100011001001110100010101000110010011101 :
(key == 11'b11110101111) ? 46'b0001010100000111001101000010101000001110011010 :
(key == 11'b11110110000) ? 46'b0001010011110101001011100010100111101010010111 :
(key == 11'b11110110001) ? 46'b0001010011100011001011000010100111000110010110 :
(key == 11'b11110110010) ? 46'b0001010011010001001100000010100110100010011000 :
(key == 11'b11110110011) ? 46'b0001010010111111001110000010100101111110011100 :
(key == 11'b11110110100) ? 46'b0001010010101101010001000010100101011010100010 :
(key == 11'b11110110101) ? 46'b0001010010011011010100000010100100110110101000 :
(key == 11'b11110110110) ? 46'b0001010010001001011000000010100100010010110000 :
(key == 11'b11110110111) ? 46'b0001010001110111011101000010100011101110111010 :
(key == 11'b11110111000) ? 46'b0001010001100101100011100010100011001011000111 :
(key == 11'b11110111001) ? 46'b0001010001010011101010000010100010100111010100 :
(key == 11'b11110111010) ? 46'b0001010001000001110001100010100010000011100011 :
(key == 11'b11110111011) ? 46'b0001010000101111111010000010100001011111110100 :
(key == 11'b11110111100) ? 46'b0001010000011110000100000010100000111100001000 :
(key == 11'b11110111101) ? 46'b0001010000001100001110000010100000011000011100 :
(key == 11'b11110111110) ? 46'b0001001111111010011001000010011111110100110010 :
(key == 11'b11110111111) ? 46'b0001001111101000100101000010011111010001001010 :
(key == 11'b11111000000) ? 46'b0001001111010110110010000010011110101101100100 :
(key == 11'b11111000001) ? 46'b0001001111000101000000000010011110001010000000 :
(key == 11'b11111000010) ? 46'b0001001110110011001111000010011101100110011110 :
(key == 11'b11111000011) ? 46'b0001001110100001011110000010011101000010111100 :
(key == 11'b11111000100) ? 46'b0001001110001111101110100010011100011111011101 :
(key == 11'b11111000101) ? 46'b0001001101111110000000000010011011111100000000 :
(key == 11'b11111000110) ? 46'b0001001101101100010010000010011011011000100100 :
(key == 11'b11111000111) ? 46'b0001001101011010100100100010011010110101001001 :
(key == 11'b11111001000) ? 46'b0001001101001000111000100010011010010001110001 :
(key == 11'b11111001001) ? 46'b0001001100110111001101000010011001101110011010 :
(key == 11'b11111001010) ? 46'b0001001100100101100010000010011001001011000100 :
(key == 11'b11111001011) ? 46'b0001001100010011111000000010011000100111110000 :
(key == 11'b11111001100) ? 46'b0001001100000010010000000010011000000100100000 :
(key == 11'b11111001101) ? 46'b0001001011110000101000000010010111100001010000 :
(key == 11'b11111001110) ? 46'b0001001011011111000001000010010110111110000010 :
(key == 11'b11111001111) ? 46'b0001001011001101011010100010010110011010110101 :
(key == 11'b11111010000) ? 46'b0001001010111011110101000010010101110111101010 :
(key == 11'b11111010001) ? 46'b0001001010101010010000000010010101010100100000 :
(key == 11'b11111010010) ? 46'b0001001010011000101100100010010100110001011001 :
(key == 11'b11111010011) ? 46'b0001001010000111001010000010010100001110010100 :
(key == 11'b11111010100) ? 46'b0001001001110101100111100010010011101011001111 :
(key == 11'b11111010101) ? 46'b0001001001100100000110000010010011001000001100 :
(key == 11'b11111010110) ? 46'b0001001001010010100110000010010010100101001100 :
(key == 11'b11111010111) ? 46'b0001001001000001000110100010010010000010001101 :
(key == 11'b11111011000) ? 46'b0001001000101111101000000010010001011111010000 :
(key == 11'b11111011001) ? 46'b0001001000011110001010000010010000111100010100 :
(key == 11'b11111011010) ? 46'b0001001000001100101101000010010000011001011010 :
(key == 11'b11111011011) ? 46'b0001000111111011010001000010001111110110100010 :
(key == 11'b11111011100) ? 46'b0001000111101001110101100010001111010011101011 :
(key == 11'b11111011101) ? 46'b0001000111011000011010100010001110110000110101 :
(key == 11'b11111011110) ? 46'b0001000111000111000001000010001110001110000010 :
(key == 11'b11111011111) ? 46'b0001000110110101101000000010001101101011010000 :
(key == 11'b11111100000) ? 46'b0001000110100100001111100010001101001000011111 :
(key == 11'b11111100001) ? 46'b0001000110010010111000000010001100100101110000 :
(key == 11'b11111100010) ? 46'b0001000110000001100010000010001100000011000100 :
(key == 11'b11111100011) ? 46'b0001000101110000001101000010001011100000011010 :
(key == 11'b11111100100) ? 46'b0001000101011110111000000010001010111101110000 :
(key == 11'b11111100101) ? 46'b0001000101001101100011100010001010011011000111 :
(key == 11'b11111100110) ? 46'b0001000100111100010000000010001001111000100000 :
(key == 11'b11111100111) ? 46'b0001000100101010111110000010001001010101111100 :
(key == 11'b11111101000) ? 46'b0001000100011001101101000010001000110011011010 :
(key == 11'b11111101001) ? 46'b0001000100001000011100100010001000010000111001 :
(key == 11'b11111101010) ? 46'b0001000011110111001100100010000111101110011001 :
(key == 11'b11111101011) ? 46'b0001000011100101111101000010000111001011111010 :
(key == 11'b11111101100) ? 46'b0001000011010100101111100010000110101001011111 :
(key == 11'b11111101101) ? 46'b0001000011000011100001100010000110000111000011 :
(key == 11'b11111101110) ? 46'b0001000010110010010101100010000101100100101011 :
(key == 11'b11111101111) ? 46'b0001000010100001001001100010000101000010010011 :
(key == 11'b11111110000) ? 46'b0001000010001111111111000010000100011111111110 :
(key == 11'b11111110001) ? 46'b0001000001111110110100100010000011111101101001 :
(key == 11'b11111110010) ? 46'b0001000001101101101011000010000011011011010110 :
(key == 11'b11111110011) ? 46'b0001000001011100100010000010000010111001000100 :
(key == 11'b11111110100) ? 46'b0001000001001011011010100010000010010110110101 :
(key == 11'b11111110101) ? 46'b0001000000111010010011100010000001110100100111 :
(key == 11'b11111110110) ? 46'b0001000000101001001101100010000001010010011011 :
(key == 11'b11111110111) ? 46'b0001000000011000001000000010000000110000010000 :
(key == 11'b11111111000) ? 46'b0001000000000111000011100010000000001110000111 :
(key == 11'b11111111001) ? 46'b0000111111110110000000000001111111101100000000 :
(key == 11'b11111111010) ? 46'b0000111111100100111101000001111111001001111010 :
(key == 11'b11111111011) ? 46'b0000111111010011111011000001111110100111110110 :
(key == 11'b11111111100) ? 46'b0000111111000010111010000001111110000101110100 :
(key == 11'b11111111101) ? 46'b0000111110110001111001000001111101100011110010 :
(key == 11'b11111111110) ? 46'b0000111110100000111001100001111101000001110011 :
(key == 11'b11111111111) ? 46'b0000111110001111111010100001111100011111110101 : 46'd0;

endmodule

`default_nettype wire
