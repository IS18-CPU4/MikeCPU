`default_nettype none

module finv
   ( input wire [31:0] x,
     output wire [31:0] y,
     output wire ovf);

   /* TODO: assumptions
    * - inputs and output are not unnormal numbers or NaN or +-inf 
    * - if e is 0, the number is interpreted as +0
    * - overflow and underflow are treated as the same for ovf wire
    * - when underflow, y will be 0
    */

   // split sequence to each subsequence
   wire xs;
   wire [7:0] xe;
   wire [22:0] xm;
   assign {xs, xe, xm} = x;

   // calc s
   wire s;
   assign s = xs;

   // calc e
   wire [7:0] e;
   assign e = (xm == 23'd0) ? 8'd254 - xe : 8'd253 - xe; 

   // calc m
   wire [22:0] m;
   wire [45:0] val;
   wire [10:0] key;
   wire [11:0] v;
   assign {key, v} = xm;
   // lookup table and get constant and grad
   lookup_table lt(key, val);
   wire [24:0] constant;
   wire [22:0] grad;
   // constant supplements 1 at the MSB
   assign constant = {1'b1, val[45:23], 1'b0};
   assign grad = val[22:0];
   wire [46:0] grad2; // length 47 = 24 + 23
   assign grad2 = {1'b1, xm, 1'b0} * grad;
   wire [23:0] tmp_m;
   assign tmp_m = constant - grad2[46:23];
   // assign tmp_m = constant - {1'b0, grad2[46:24]};
   assign m = (xm == 23'd0) ? 23'd0 : {tmp_m[21:0], 1'b0};

   assign y = {s, e, m};
   assign ovf = 0;

endmodule

module lookup_table
   ( input wire [10:0] key,
     output wire [45:0] value);

   assign value =
(key == 11'b00000000000) ? 46'b1111111111100000000000111111111111000000000001 :
(key == 11'b00000000001) ? 46'b1111111110100000000100111111111101000000001101 :
(key == 11'b00000000010) ? 46'b1111111101100000001100111111111011000000100101 :
(key == 11'b00000000011) ? 46'b1111111100100000011000111111111001000001001001 :
(key == 11'b00000000100) ? 46'b1111111011100000101000111111110111000001111001 :
(key == 11'b00000000101) ? 46'b1111111010100000111100111111110101000010110101 :
(key == 11'b00000000110) ? 46'b1111111001100001010100011111110011000011111100 :
(key == 11'b00000000111) ? 46'b1111111000100001110000011111110001000101001111 :
(key == 11'b00000001000) ? 46'b1111110111100010010000011111101111000110101111 :
(key == 11'b00000001001) ? 46'b1111110110100010110011111111101101001000011010 :
(key == 11'b00000001010) ? 46'b1111110101100011011011111111101011001010010001 :
(key == 11'b00000001011) ? 46'b1111110100100100000111011111101001001100010011 :
(key == 11'b00000001100) ? 46'b1111110011100100110110111111100111001110100001 :
(key == 11'b00000001101) ? 46'b1111110010100101101010011111100101010000111011 :
(key == 11'b00000001110) ? 46'b1111110001100110100001111111100011010011100001 :
(key == 11'b00000001111) ? 46'b1111110000100111011101011111100001010110010011 :
(key == 11'b00000010000) ? 46'b1111101111101000011100011111011111011001010000 :
(key == 11'b00000010001) ? 46'b1111101110101001011111111111011101011100011001 :
(key == 11'b00000010010) ? 46'b1111101101101010100110111111011011011111101101 :
(key == 11'b00000010011) ? 46'b1111101100101011110001111111011001100011001101 :
(key == 11'b00000010100) ? 46'b1111101011101101000000011111010111100110111000 :
(key == 11'b00000010101) ? 46'b1111101010101110010011011111010101101010101111 :
(key == 11'b00000010110) ? 46'b1111101001101111101001111111010011101110110001 :
(key == 11'b00000010111) ? 46'b1111101000110001000100011111010001110010111111 :
(key == 11'b00000011000) ? 46'b1111100111110010100010111111001111110111011001 :
(key == 11'b00000011001) ? 46'b1111100110110100000100111111001101111011111101 :
(key == 11'b00000011010) ? 46'b1111100101110101101010111111001100000000101110 :
(key == 11'b00000011011) ? 46'b1111100100110111010100111111001010000101101001 :
(key == 11'b00000011100) ? 46'b1111100011111001000010011111001000001010110000 :
(key == 11'b00000011101) ? 46'b1111100010111010110100011111000110010000000011 :
(key == 11'b00000011110) ? 46'b1111100001111100101001011111000100010101100000 :
(key == 11'b00000011111) ? 46'b1111100000111110100010111111000010011011001010 :
(key == 11'b00000100000) ? 46'b1111100000000000011111111111000000100000111110 :
(key == 11'b00000100001) ? 46'b1111011111000010100000111110111110100110111110 :
(key == 11'b00000100010) ? 46'b1111011110000100100101011110111100101101001000 :
(key == 11'b00000100011) ? 46'b1111011101000110101101111110111010110011011110 :
(key == 11'b00000100100) ? 46'b1111011100001000111010011110111000111010000000 :
(key == 11'b00000100101) ? 46'b1111011011001011001010011110110111000000101100 :
(key == 11'b00000100110) ? 46'b1111011010001101011110011110110101000111100100 :
(key == 11'b00000100111) ? 46'b1111011001001111110101111110110011001110100110 :
(key == 11'b00000101000) ? 46'b1111011000010010010001011110110001010101110100 :
(key == 11'b00000101001) ? 46'b1111010111010100110000011110101111011101001101 :
(key == 11'b00000101010) ? 46'b1111010110010111010011011110101101100100110001 :
(key == 11'b00000101011) ? 46'b1111010101011001111010011110101011101100100000 :
(key == 11'b00000101100) ? 46'b1111010100011100100100111110101001110100011011 :
(key == 11'b00000101101) ? 46'b1111010011011111010010111110100111111100011111 :
(key == 11'b00000101110) ? 46'b1111010010100010000100111110100110000100101111 :
(key == 11'b00000101111) ? 46'b1111010001100100111010011110100100001101001010 :
(key == 11'b00000110000) ? 46'b1111010000100111110011111110100010010101110000 :
(key == 11'b00000110001) ? 46'b1111001111101010110001011110100000011110100010 :
(key == 11'b00000110010) ? 46'b1111001110101101110010011110011110100111011110 :
(key == 11'b00000110011) ? 46'b1111001101110000110110111110011100110000100100 :
(key == 11'b00000110100) ? 46'b1111001100110011111110111110011010111001110101 :
(key == 11'b00000110101) ? 46'b1111001011110111001011011110011001000011010010 :
(key == 11'b00000110110) ? 46'b1111001010111010011010111110010111001100111001 :
(key == 11'b00000110111) ? 46'b1111001001111101101110011110010101010110101011 :
(key == 11'b00000111000) ? 46'b1111001001000001000101011110010011100000101000 :
(key == 11'b00000111001) ? 46'b1111001000000100100000011110010001101010110000 :
(key == 11'b00000111010) ? 46'b1111000111000111111110111110001111110101000010 :
(key == 11'b00000111011) ? 46'b1111000110001011100000111110001101111111011111 :
(key == 11'b00000111100) ? 46'b1111000101001111000110111110001100001010000111 :
(key == 11'b00000111101) ? 46'b1111000100010010110000011110001010010100111010 :
(key == 11'b00000111110) ? 46'b1111000011010110011101011110001000011111110110 :
(key == 11'b00000111111) ? 46'b1111000010011010001110011110000110101010111110 :
(key == 11'b00001000000) ? 46'b1111000001011110000010111110000100110110010001 :
(key == 11'b00001000001) ? 46'b1111000000100001111010111110000011000001101110 :
(key == 11'b00001000010) ? 46'b1110111111100101110110111110000001001101010110 :
(key == 11'b00001000011) ? 46'b1110111110101001110101111101111111011001000111 :
(key == 11'b00001000100) ? 46'b1110111101101101111001011101111101100101000101 :
(key == 11'b00001000101) ? 46'b1110111100110001111111111101111011110001001100 :
(key == 11'b00001000110) ? 46'b1110111011110110001001111101111001111101011101 :
(key == 11'b00001000111) ? 46'b1110111010111010010111111101111000001001111001 :
(key == 11'b00001001000) ? 46'b1110111001111110101001011101110110010110100000 :
(key == 11'b00001001001) ? 46'b1110111001000010111110011101110100100011010001 :
(key == 11'b00001001010) ? 46'b1110111000000111010111011101110010110000001101 :
(key == 11'b00001001011) ? 46'b1110110111001011110011011101110000111101010010 :
(key == 11'b00001001100) ? 46'b1110110110010000010011011101101111001010100011 :
(key == 11'b00001001101) ? 46'b1110110101010100110110111101101101010111111101 :
(key == 11'b00001001110) ? 46'b1110110100011001011101111101101011100101100010 :
(key == 11'b00001001111) ? 46'b1110110011011110001000011101101001110011010001 :
(key == 11'b00001010000) ? 46'b1110110010100010110110111101101000000001001011 :
(key == 11'b00001010001) ? 46'b1110110001100111101000011101100110001111001111 :
(key == 11'b00001010010) ? 46'b1110110000101100011101111101100100011101011101 :
(key == 11'b00001010011) ? 46'b1110101111110001010110011101100010101011110101 :
(key == 11'b00001010100) ? 46'b1110101110110110010010111101100000111010011000 :
(key == 11'b00001010101) ? 46'b1110101101111011010010111101011111001001000101 :
(key == 11'b00001010110) ? 46'b1110101101000000010110011101011101010111111100 :
(key == 11'b00001010111) ? 46'b1110101100000101011101011101011011100110111101 :
(key == 11'b00001011000) ? 46'b1110101011001010100111111101011001110110001000 :
(key == 11'b00001011001) ? 46'b1110101010001111110101111101011000000101011110 :
(key == 11'b00001011010) ? 46'b1110101001010101000111111101010110010100111110 :
(key == 11'b00001011011) ? 46'b1110101000011010011100111101010100100100101000 :
(key == 11'b00001011100) ? 46'b1110100111011111110101011101010010110100011011 :
(key == 11'b00001011101) ? 46'b1110100110100101010001011101010001000100011001 :
(key == 11'b00001011110) ? 46'b1110100101101010110000111101001111010100100000 :
(key == 11'b00001011111) ? 46'b1110100100110000010100011101001101100100110011 :
(key == 11'b00001100000) ? 46'b1110100011110101111010111101001011110101001111 :
(key == 11'b00001100001) ? 46'b1110100010111011100100111101001010000101110101 :
(key == 11'b00001100010) ? 46'b1110100010000001010010011101001000010110100100 :
(key == 11'b00001100011) ? 46'b1110100001000111000011011101000110100111011110 :
(key == 11'b00001100100) ? 46'b1110100000001100110111111101000100111000100010 :
(key == 11'b00001100101) ? 46'b1110011111010010101111111101000011001001101111 :
(key == 11'b00001100110) ? 46'b1110011110011000101011011101000001011011000111 :
(key == 11'b00001100111) ? 46'b1110011101011110101010011100111111101100101001 :
(key == 11'b00001101000) ? 46'b1110011100100100101100011100111101111110010011 :
(key == 11'b00001101001) ? 46'b1110011011101010110010011100111100010000001001 :
(key == 11'b00001101010) ? 46'b1110011010110000111011011100111010100010000111 :
(key == 11'b00001101011) ? 46'b1110011001110111001000011100111000110100010000 :
(key == 11'b00001101100) ? 46'b1110011000111101011000011100110111000110100011 :
(key == 11'b00001101101) ? 46'b1110011000000011101011111100110101011000111111 :
(key == 11'b00001101110) ? 46'b1110010111001010000010111100110011101011100101 :
(key == 11'b00001101111) ? 46'b1110010110010000011100111100110001111110010100 :
(key == 11'b00001110000) ? 46'b1110010101010110111010111100110000010001001110 :
(key == 11'b00001110001) ? 46'b1110010100011101011011111100101110100100010001 :
(key == 11'b00001110010) ? 46'b1110010011100100000000011100101100110111011101 :
(key == 11'b00001110011) ? 46'b1110010010101010101000011100101011001010110100 :
(key == 11'b00001110100) ? 46'b1110010001110001010011111100101001011110010100 :
(key == 11'b00001110101) ? 46'b1110010000111000000010011100100111110001111101 :
(key == 11'b00001110110) ? 46'b1110001111111110110100111100100110000101110001 :
(key == 11'b00001110111) ? 46'b1110001111000101101010011100100100011001101110 :
(key == 11'b00001111000) ? 46'b1110001110001100100011011100100010101101110100 :
(key == 11'b00001111001) ? 46'b1110001101010011011111011100100001000010000100 :
(key == 11'b00001111010) ? 46'b1110001100011010011110111100011111010110011101 :
(key == 11'b00001111011) ? 46'b1110001011100001100001111100011101101011000000 :
(key == 11'b00001111100) ? 46'b1110001010101000101000011100011011111111101101 :
(key == 11'b00001111101) ? 46'b1110001001101111110001111100011010010100100011 :
(key == 11'b00001111110) ? 46'b1110001000110110111110111100011000101001100010 :
(key == 11'b00001111111) ? 46'b1110000111111110001111011100010110111110101011 :
(key == 11'b00010000000) ? 46'b1110000111000101100010111100010101010011111101 :
(key == 11'b00010000001) ? 46'b1110000110001100111010011100010011101001011001 :
(key == 11'b00010000010) ? 46'b1110000101010100010100011100010001111110111110 :
(key == 11'b00010000011) ? 46'b1110000100011011110010011100010000010100101101 :
(key == 11'b00010000100) ? 46'b1110000011100011010011011100001110101010100101 :
(key == 11'b00010000101) ? 46'b1110000010101010110111011100001101000000100101 :
(key == 11'b00010000110) ? 46'b1110000001110010011111011100001011010110110000 :
(key == 11'b00010000111) ? 46'b1110000000111010001010011100001001101101000100 :
(key == 11'b00010001000) ? 46'b1110000000000001111000011100001000000011100001 :
(key == 11'b00010001001) ? 46'b1101111111001001101001111100000110011010000111 :
(key == 11'b00010001010) ? 46'b1101111110010001011110111100000100110000110111 :
(key == 11'b00010001011) ? 46'b1101111101011001010110111100000011000111101111 :
(key == 11'b00010001100) ? 46'b1101111100100001010010011100000001011110110010 :
(key == 11'b00010001101) ? 46'b1101111011101001010000111011111111110101111101 :
(key == 11'b00010001110) ? 46'b1101111010110001010010111011111110001101010001 :
(key == 11'b00010001111) ? 46'b1101111001111001010111111011111100100100101110 :
(key == 11'b00010010000) ? 46'b1101111001000001100000011011111010111100010101 :
(key == 11'b00010010001) ? 46'b1101111000001001101100011011111001010100000101 :
(key == 11'b00010010010) ? 46'b1101110111010001111011011011110111101011111110 :
(key == 11'b00010010011) ? 46'b1101110110011010001101011011110110000100000000 :
(key == 11'b00010010100) ? 46'b1101110101100010100010111011110100011100001011 :
(key == 11'b00010010101) ? 46'b1101110100101010111011111011110010110100100000 :
(key == 11'b00010010110) ? 46'b1101110011110011010111111011110001001100111101 :
(key == 11'b00010010111) ? 46'b1101110010111011110110111011101111100101100011 :
(key == 11'b00010011000) ? 46'b1101110010000100011001011011101101111110010011 :
(key == 11'b00010011001) ? 46'b1101110001001100111110111011101100010111001011 :
(key == 11'b00010011010) ? 46'b1101110000010101100111111011101010110000001100 :
(key == 11'b00010011011) ? 46'b1101101111011110010011111011101001001001010111 :
(key == 11'b00010011100) ? 46'b1101101110100111000011011011100111100010101010 :
(key == 11'b00010011101) ? 46'b1101101101101111110101111011100101111100000110 :
(key == 11'b00010011110) ? 46'b1101101100111000101011111011100100010101101100 :
(key == 11'b00010011111) ? 46'b1101101100000001100100011011100010101111011001 :
(key == 11'b00010100000) ? 46'b1101101011001010100000111011100001001001010001 :
(key == 11'b00010100001) ? 46'b1101101010010011011111111011011111100011010000 :
(key == 11'b00010100010) ? 46'b1101101001011100100010011011011101111101011001 :
(key == 11'b00010100011) ? 46'b1101101000100101101000011011011100010111101011 :
(key == 11'b00010100100) ? 46'b1101100111101110110000111011011010110010000101 :
(key == 11'b00010100101) ? 46'b1101100110110111111100111011011001001100101000 :
(key == 11'b00010100110) ? 46'b1101100110000001001100011011010111100111010100 :
(key == 11'b00010100111) ? 46'b1101100101001010011110011011010110000010001000 :
(key == 11'b00010101000) ? 46'b1101100100010011110011111011010100011101000110 :
(key == 11'b00010101001) ? 46'b1101100011011101001100111011010010111000001101 :
(key == 11'b00010101010) ? 46'b1101100010100110101000011011010001010011011011 :
(key == 11'b00010101011) ? 46'b1101100001110000000111011011001111101110110011 :
(key == 11'b00010101100) ? 46'b1101100000111001101001111011001110001010010100 :
(key == 11'b00010101101) ? 46'b1101100000000011001110111011001100100101111100 :
(key == 11'b00010101110) ? 46'b1101011111001100110111011011001011000001101110 :
(key == 11'b00010101111) ? 46'b1101011110010110100010111011001001011101101001 :
(key == 11'b00010110000) ? 46'b1101011101100000010001011011000111111001101100 :
(key == 11'b00010110001) ? 46'b1101011100101010000011011011000110010101111000 :
(key == 11'b00010110010) ? 46'b1101011011110011110111111011000100110010001011 :
(key == 11'b00010110011) ? 46'b1101011010111101101111111011000011001110101000 :
(key == 11'b00010110100) ? 46'b1101011010000111101010111011000001101011001101 :
(key == 11'b00010110101) ? 46'b1101011001010001101001011011000000000111111100 :
(key == 11'b00010110110) ? 46'b1101011000011011101010111010111110100100110011 :
(key == 11'b00010110111) ? 46'b1101010111100101101110111010111101000001110001 :
(key == 11'b00010111000) ? 46'b1101010110101111110110011010111011011110111001 :
(key == 11'b00010111001) ? 46'b1101010101111010000000111010111001111100001000 :
(key == 11'b00010111010) ? 46'b1101010101000100001110111010111000011001100010 :
(key == 11'b00010111011) ? 46'b1101010100001110011111011010110110110111000010 :
(key == 11'b00010111100) ? 46'b1101010011011000110011011010110101010100101100 :
(key == 11'b00010111101) ? 46'b1101010010100011001010011010110011110010011110 :
(key == 11'b00010111110) ? 46'b1101010001101101100100011010110010010000011000 :
(key == 11'b00010111111) ? 46'b1101010000111000000001011010110000101110011011 :
(key == 11'b00011000000) ? 46'b1101010000000010100001011010101111001100100110 :
(key == 11'b00011000001) ? 46'b1101001111001101000100011010101101101010111001 :
(key == 11'b00011000010) ? 46'b1101001110010111101010011010101100001001010101 :
(key == 11'b00011000011) ? 46'b1101001101100010010011111010101010100111111010 :
(key == 11'b00011000100) ? 46'b1101001100101100111111111010101001000110100110 :
(key == 11'b00011000101) ? 46'b1101001011110111101111011010100111100101011011 :
(key == 11'b00011000110) ? 46'b1101001011000010100001111010100110000100011000 :
(key == 11'b00011000111) ? 46'b1101001010001101010110111010100100100011011101 :
(key == 11'b00011001000) ? 46'b1101001001011000001111011010100011000010101011 :
(key == 11'b00011001001) ? 46'b1101001000100011001010111010100001100010000001 :
(key == 11'b00011001010) ? 46'b1101000111101110001001011010100000000001011111 :
(key == 11'b00011001011) ? 46'b1101000110111001001010111010011110100001000110 :
(key == 11'b00011001100) ? 46'b1101000110000100001111011010011101000000110101 :
(key == 11'b00011001101) ? 46'b1101000101001111010110111010011011100000101011 :
(key == 11'b00011001110) ? 46'b1101000100011010100001011010011010000000101011 :
(key == 11'b00011001111) ? 46'b1101000011100101101110111010011000100000110010 :
(key == 11'b00011010000) ? 46'b1101000010110000111111011010010111000001000001 :
(key == 11'b00011010001) ? 46'b1101000001111100010010111010010101100001011001 :
(key == 11'b00011010010) ? 46'b1101000001000111101001011010010100000001111001 :
(key == 11'b00011010011) ? 46'b1101000000010011000010011010010010100010100000 :
(key == 11'b00011010100) ? 46'b1100111111011110011110111010010001000011010000 :
(key == 11'b00011010101) ? 46'b1100111110101001111110011010001111100100001000 :
(key == 11'b00011010110) ? 46'b1100111101110101100000111010001110000101001000 :
(key == 11'b00011010111) ? 46'b1100111101000001000101111010001100100110010000 :
(key == 11'b00011011000) ? 46'b1100111100001100101110011010001011000111100000 :
(key == 11'b00011011001) ? 46'b1100111011011000011001011010001001101000111000 :
(key == 11'b00011011010) ? 46'b1100111010100100000111111010001000001010011000 :
(key == 11'b00011011011) ? 46'b1100111001101111111000111010000110101100000000 :
(key == 11'b00011011100) ? 46'b1100111000111011101100111010000101001101110000 :
(key == 11'b00011011101) ? 46'b1100111000000111100011111010000011101111101000 :
(key == 11'b00011011110) ? 46'b1100110111010011011101111010000010010001101000 :
(key == 11'b00011011111) ? 46'b1100110110011111011010111010000000110011110001 :
(key == 11'b00011100000) ? 46'b1100110101101011011010111001111111010110000001 :
(key == 11'b00011100001) ? 46'b1100110100110111011101011001111101111000011000 :
(key == 11'b00011100010) ? 46'b1100110100000011100011011001111100011010111001 :
(key == 11'b00011100011) ? 46'b1100110011001111101011111001111010111101100000 :
(key == 11'b00011100100) ? 46'b1100110010011011110111011001111001100000001111 :
(key == 11'b00011100101) ? 46'b1100110001101000000101111001111000000011000111 :
(key == 11'b00011100110) ? 46'b1100110000110100010111011001110110100110000110 :
(key == 11'b00011100111) ? 46'b1100110000000000101011011001110101001001001101 :
(key == 11'b00011101000) ? 46'b1100101111001101000010111001110011101100011101 :
(key == 11'b00011101001) ? 46'b1100101110011001011100111001110010001111110011 :
(key == 11'b00011101010) ? 46'b1100101101100101111001111001110000110011010010 :
(key == 11'b00011101011) ? 46'b1100101100110010011001011001101111010110110111 :
(key == 11'b00011101100) ? 46'b1100101011111110111100011001101101111010100110 :
(key == 11'b00011101101) ? 46'b1100101011001011100001111001101100011110011011 :
(key == 11'b00011101110) ? 46'b1100101010011000001010011001101011000010011001 :
(key == 11'b00011101111) ? 46'b1100101001100100110101111001101001100110011110 :
(key == 11'b00011110000) ? 46'b1100101000110001100011111001101000001010101011 :
(key == 11'b00011110001) ? 46'b1100100111111110010100111001100110101110111111 :
(key == 11'b00011110010) ? 46'b1100100111001011001000111001100101010011011100 :
(key == 11'b00011110011) ? 46'b1100100110010111111111111001100011111000000000 :
(key == 11'b00011110100) ? 46'b1100100101100100111001011001100010011100101011 :
(key == 11'b00011110101) ? 46'b1100100100110001110101111001100001000001011111 :
(key == 11'b00011110110) ? 46'b1100100011111110110101011001011111100110011010 :
(key == 11'b00011110111) ? 46'b1100100011001011110111011001011110001011011100 :
(key == 11'b00011111000) ? 46'b1100100010011000111100111001011100110000100111 :
(key == 11'b00011111001) ? 46'b1100100001100110000100011001011011010101111000 :
(key == 11'b00011111010) ? 46'b1100100000110011001111011001011001111011010010 :
(key == 11'b00011111011) ? 46'b1100100000000000011100111001011000100000110011 :
(key == 11'b00011111100) ? 46'b1100011111001101101101011001010111000110011011 :
(key == 11'b00011111101) ? 46'b1100011110011011000000011001010101101100001011 :
(key == 11'b00011111110) ? 46'b1100011101101000010110011001010100010010000010 :
(key == 11'b00011111111) ? 46'b1100011100110101101111011001010010111000000001 :
(key == 11'b00100000000) ? 46'b1100011100000011001010111001010001011110001000 :
(key == 11'b00100000001) ? 46'b1100011011010000101001011001010000000100010110 :
(key == 11'b00100000010) ? 46'b1100011010011110001010111001001110101010101100 :
(key == 11'b00100000011) ? 46'b1100011001101011101110111001001101010001001000 :
(key == 11'b00100000100) ? 46'b1100011000111001010101111001001011110111101101 :
(key == 11'b00100000101) ? 46'b1100011000000110111111011001001010011110011001 :
(key == 11'b00100000110) ? 46'b1100010111010100101011111001001001000101001100 :
(key == 11'b00100000111) ? 46'b1100010110100010011010111001000111101100000110 :
(key == 11'b00100001000) ? 46'b1100010101110000001100111001000110010011001000 :
(key == 11'b00100001001) ? 46'b1100010100111110000001111001000100111010010010 :
(key == 11'b00100001010) ? 46'b1100010100001011111001011001000011100001100010 :
(key == 11'b00100001011) ? 46'b1100010011011001110011111001000010001000111011 :
(key == 11'b00100001100) ? 46'b1100010010100111110000111001000000110000011010 :
(key == 11'b00100001101) ? 46'b1100010001110101110000111000111111011000000001 :
(key == 11'b00100001110) ? 46'b1100010001000011110011011000111101111111101111 :
(key == 11'b00100001111) ? 46'b1100010000010001111000111000111100100111100101 :
(key == 11'b00100010000) ? 46'b1100001111100000000000111000111011001111100001 :
(key == 11'b00100010001) ? 46'b1100001110101110001011111000111001110111100101 :
(key == 11'b00100010010) ? 46'b1100001101111100011001011000111000011111110000 :
(key == 11'b00100010011) ? 46'b1100001101001010101001111000110111001000000011 :
(key == 11'b00100010100) ? 46'b1100001100011000111100111000110101110000011101 :
(key == 11'b00100010101) ? 46'b1100001011100111010010111000110100011000111110 :
(key == 11'b00100010110) ? 46'b1100001010110101101011011000110011000001100110 :
(key == 11'b00100010111) ? 46'b1100001010000100000110011000110001101010010101 :
(key == 11'b00100011000) ? 46'b1100001001010010100100111000110000010011001100 :
(key == 11'b00100011001) ? 46'b1100001000100001000101011000101110111100001010 :
(key == 11'b00100011010) ? 46'b1100000111101111101000111000101101100101001111 :
(key == 11'b00100011011) ? 46'b1100000110111110001110111000101100001110011010 :
(key == 11'b00100011100) ? 46'b1100000110001100110111111000101010110111101110 :
(key == 11'b00100011101) ? 46'b1100000101011011100011011000101001100001001000 :
(key == 11'b00100011110) ? 46'b1100000100101010010001111000101000001010101010 :
(key == 11'b00100011111) ? 46'b1100000011111001000010111000100110110100010010 :
(key == 11'b00100100000) ? 46'b1100000011000111110110011000100101011110000010 :
(key == 11'b00100100001) ? 46'b1100000010010110101100111000100100000111111001 :
(key == 11'b00100100010) ? 46'b1100000001100101100110011000100010110001110111 :
(key == 11'b00100100011) ? 46'b1100000000110100100001111000100001011011111100 :
(key == 11'b00100100100) ? 46'b1100000000000011100000011000100000000110001000 :
(key == 11'b00100100101) ? 46'b1011111111010010100001011000011110110000011011 :
(key == 11'b00100100110) ? 46'b1011111110100001100101011000011101011010110101 :
(key == 11'b00100100111) ? 46'b1011111101110000101011111000011100000101010110 :
(key == 11'b00100101000) ? 46'b1011111100111111110100111000011010101111111110 :
(key == 11'b00100101001) ? 46'b1011111100001111000000111000011001011010101101 :
(key == 11'b00100101010) ? 46'b1011111011011110001111011000011000000101100011 :
(key == 11'b00100101011) ? 46'b1011111010101101100000011000010110110000100000 :
(key == 11'b00100101100) ? 46'b1011111001111100110100011000010101011011100100 :
(key == 11'b00100101101) ? 46'b1011111001001100001010111000010100000110101111 :
(key == 11'b00100101110) ? 46'b1011111000011011100011111000010010110010000000 :
(key == 11'b00100101111) ? 46'b1011110111101010111111111000010001011101011010 :
(key == 11'b00100110000) ? 46'b1011110110111010011101111000010000001000111001 :
(key == 11'b00100110001) ? 46'b1011110110001001111110111000001110110100011111 :
(key == 11'b00100110010) ? 46'b1011110101011001100010111000001101100000001101 :
(key == 11'b00100110011) ? 46'b1011110100101001001000111000001100001100000001 :
(key == 11'b00100110100) ? 46'b1011110011111000110001111000001010110111111100 :
(key == 11'b00100110101) ? 46'b1011110011001000011101011000001001100011111110 :
(key == 11'b00100110110) ? 46'b1011110010011000001011111000001000010000000111 :
(key == 11'b00100110111) ? 46'b1011110001100111111100011000000110111100010110 :
(key == 11'b00100111000) ? 46'b1011110000110111101111111000000101101000101101 :
(key == 11'b00100111001) ? 46'b1011110000000111100101111000000100010101001010 :
(key == 11'b00100111010) ? 46'b1011101111010111011110111000000011000001101110 :
(key == 11'b00100111011) ? 46'b1011101110100111011001111000000001101110011001 :
(key == 11'b00100111100) ? 46'b1011101101110111010111111000000000011011001011 :
(key == 11'b00100111101) ? 46'b1011101101000111011000010111111111001000000011 :
(key == 11'b00100111110) ? 46'b1011101100010111011011010111111101110101000010 :
(key == 11'b00100111111) ? 46'b1011101011100111100000110111111100100010001000 :
(key == 11'b00101000000) ? 46'b1011101010110111101001010111111011001111010101 :
(key == 11'b00101000001) ? 46'b1011101010000111110011110111111001111100100111 :
(key == 11'b00101000010) ? 46'b1011101001011000000001010111111000101010000001 :
(key == 11'b00101000011) ? 46'b1011101000101000010001010111110111010111100010 :
(key == 11'b00101000100) ? 46'b1011100111111000100011110111110110000101001001 :
(key == 11'b00101000101) ? 46'b1011100111001000111000110111110100110010110111 :
(key == 11'b00101000110) ? 46'b1011100110011001010000110111110011100000101100 :
(key == 11'b00101000111) ? 46'b1011100101101001101010110111110010001110100111 :
(key == 11'b00101001000) ? 46'b1011100100111010000111110111110000111100101001 :
(key == 11'b00101001001) ? 46'b1011100100001010100111010111101111101010110001 :
(key == 11'b00101001010) ? 46'b1011100011011011001000110111101110011001000000 :
(key == 11'b00101001011) ? 46'b1011100010101011101101010111101101000111010101 :
(key == 11'b00101001100) ? 46'b1011100001111100010100110111101011110101110011 :
(key == 11'b00101001101) ? 46'b1011100001001100111110010111101010100100010101 :
(key == 11'b00101001110) ? 46'b1011100000011101101010010111101001010010111110 :
(key == 11'b00101001111) ? 46'b1011011111101110011000110111101000000001101110 :
(key == 11'b00101010000) ? 46'b1011011110111111001010010111100110110000100101 :
(key == 11'b00101010001) ? 46'b1011011110001111111101110111100101011111100010 :
(key == 11'b00101010010) ? 46'b1011011101100000110100010111100100001110100101 :
(key == 11'b00101010011) ? 46'b1011011100110001101100110111100010111101101111 :
(key == 11'b00101010100) ? 46'b1011011100000010101000010111100001101101000000 :
(key == 11'b00101010101) ? 46'b1011011011010011100110010111100000011100010111 :
(key == 11'b00101010110) ? 46'b1011011010100100100110110111011111001011110101 :
(key == 11'b00101010111) ? 46'b1011011001110101101001010111011101111011011000 :
(key == 11'b00101011000) ? 46'b1011011001000110101110110111011100101011000011 :
(key == 11'b00101011001) ? 46'b1011011000010111110110110111011011011010110100 :
(key == 11'b00101011010) ? 46'b1011010111101001000001010111011010001010101011 :
(key == 11'b00101011011) ? 46'b1011010110111010001110010111011000111010101001 :
(key == 11'b00101011100) ? 46'b1011010110001011011101010111010111101010101100 :
(key == 11'b00101011101) ? 46'b1011010101011100101111010111010110011010110111 :
(key == 11'b00101011110) ? 46'b1011010100101110000011110111010101001011001000 :
(key == 11'b00101011111) ? 46'b1011010011111111011010110111010011111011100000 :
(key == 11'b00101100000) ? 46'b1011010011010000110100010111010010101011111110 :
(key == 11'b00101100001) ? 46'b1011010010100010001111110111010001011100100001 :
(key == 11'b00101100010) ? 46'b1011010001110011101110010111010000001101001100 :
(key == 11'b00101100011) ? 46'b1011010001000101001111010111001110111101111101 :
(key == 11'b00101100100) ? 46'b1011010000010110110010010111001101101110110011 :
(key == 11'b00101100101) ? 46'b1011001111101000011000010111001100011111110001 :
(key == 11'b00101100110) ? 46'b1011001110111010000000010111001011010000110100 :
(key == 11'b00101100111) ? 46'b1011001110001011101011010111001010000001111111 :
(key == 11'b00101101000) ? 46'b1011001101011101011000010111001000110011001111 :
(key == 11'b00101101001) ? 46'b1011001100101111000111110111000111100100100101 :
(key == 11'b00101101010) ? 46'b1011001100000000111010010111000110010110000010 :
(key == 11'b00101101011) ? 46'b1011001011010010101110110111000101000111100101 :
(key == 11'b00101101100) ? 46'b1011001010100100100101110111000011111001001111 :
(key == 11'b00101101101) ? 46'b1011001001110110011110110111000010101010111101 :
(key == 11'b00101101110) ? 46'b1011001001001000011010110111000001011100110011 :
(key == 11'b00101101111) ? 46'b1011001000011010011001010111000000001110101111 :
(key == 11'b00101110000) ? 46'b1011000111101100011001110110111111000000110001 :
(key == 11'b00101110001) ? 46'b1011000110111110011101010110111101110010111010 :
(key == 11'b00101110010) ? 46'b1011000110010000100010110110111100100101001000 :
(key == 11'b00101110011) ? 46'b1011000101100010101010110110111011010111011101 :
(key == 11'b00101110100) ? 46'b1011000100110100110101010110111010001001111000 :
(key == 11'b00101110101) ? 46'b1011000100000111000010010110111000111100011001 :
(key == 11'b00101110110) ? 46'b1011000011011001010001110110110111101111000000 :
(key == 11'b00101110111) ? 46'b1011000010101011100011010110110110100001101101 :
(key == 11'b00101111000) ? 46'b1011000001111101110111010110110101010100100000 :
(key == 11'b00101111001) ? 46'b1011000001010000001101110110110100000111011010 :
(key == 11'b00101111010) ? 46'b1011000000100010100110110110110010111010011001 :
(key == 11'b00101111011) ? 46'b1010111111110101000010010110110001101101011111 :
(key == 11'b00101111100) ? 46'b1010111111000111100000010110110000100000101011 :
(key == 11'b00101111101) ? 46'b1010111110011010000000010110101111010011111101 :
(key == 11'b00101111110) ? 46'b1010111101101100100010110110101110000111010101 :
(key == 11'b00101111111) ? 46'b1010111100111111000111110110101100111010110011 :
(key == 11'b00110000000) ? 46'b1010111100010001101111010110101011101110010111 :
(key == 11'b00110000001) ? 46'b1010111011100100011000110110101010100010000000 :
(key == 11'b00110000010) ? 46'b1010111010110111000101010110101001010101110001 :
(key == 11'b00110000011) ? 46'b1010111010001001110011110110101000001001100111 :
(key == 11'b00110000100) ? 46'b1010111001011100100100010110100110111101100010 :
(key == 11'b00110000101) ? 46'b1010111000101111010111110110100101110001100101 :
(key == 11'b00110000110) ? 46'b1010111000000010001101010110100100100101101101 :
(key == 11'b00110000111) ? 46'b1010110111010101000101010110100011011001111011 :
(key == 11'b00110001000) ? 46'b1010110110100111111111110110100010001110001111 :
(key == 11'b00110001001) ? 46'b1010110101111010111100010110100001000010101000 :
(key == 11'b00110001010) ? 46'b1010110101001101111011110110011111110111001001 :
(key == 11'b00110001011) ? 46'b1010110100100000111101010110011110101011101111 :
(key == 11'b00110001100) ? 46'b1010110011110100000000110110011101100000011010 :
(key == 11'b00110001101) ? 46'b1010110011000111000110110110011100010101001011 :
(key == 11'b00110001110) ? 46'b1010110010011010001111110110011011001010000011 :
(key == 11'b00110001111) ? 46'b1010110001101101011010010110011001111111000000 :
(key == 11'b00110010000) ? 46'b1010110001000000100111110110011000110100000100 :
(key == 11'b00110010001) ? 46'b1010110000010011110111010110010111101001001101 :
(key == 11'b00110010010) ? 46'b1010101111100111001000110110010110011110011011 :
(key == 11'b00110010011) ? 46'b1010101110111010011101010110010101010011110001 :
(key == 11'b00110010100) ? 46'b1010101110001101110011110110010100001001001011 :
(key == 11'b00110010101) ? 46'b1010101101100001001100110110010010111110101100 :
(key == 11'b00110010110) ? 46'b1010101100110100100111110110010001110100010010 :
(key == 11'b00110010111) ? 46'b1010101100001000000101010110010000101001111110 :
(key == 11'b00110011000) ? 46'b1010101011011011100101010110001111011111110000 :
(key == 11'b00110011001) ? 46'b1010101010101111000111010110001110010101101000 :
(key == 11'b00110011010) ? 46'b1010101010000010101011110110001101001011100101 :
(key == 11'b00110011011) ? 46'b1010101001010110010010110110001100000001101001 :
(key == 11'b00110011100) ? 46'b1010101000101001111011110110001010110111110010 :
(key == 11'b00110011101) ? 46'b1010100111111101100111010110001001101110000001 :
(key == 11'b00110011110) ? 46'b1010100111010001010100110110001000100100010101 :
(key == 11'b00110011111) ? 46'b1010100110100101000100110110000111011010110000 :
(key == 11'b00110100000) ? 46'b1010100101111000110111010110000110010001010000 :
(key == 11'b00110100001) ? 46'b1010100101001100101011110110000101000111110110 :
(key == 11'b00110100010) ? 46'b1010100100100000100010110110000011111110100010 :
(key == 11'b00110100011) ? 46'b1010100011110100011011110110000010110101010010 :
(key == 11'b00110100100) ? 46'b1010100011001000010111010110000001101100001001 :
(key == 11'b00110100101) ? 46'b1010100010011100010101010110000000100011000110 :
(key == 11'b00110100110) ? 46'b1010100001110000010101010101111111011010001001 :
(key == 11'b00110100111) ? 46'b1010100001000100010111110101111110010001010001 :
(key == 11'b00110101000) ? 46'b1010100000011000011100010101111101001000011110 :
(key == 11'b00110101001) ? 46'b1010011111101100100010110101111011111111110001 :
(key == 11'b00110101010) ? 46'b1010011111000000101100010101111010110111001011 :
(key == 11'b00110101011) ? 46'b1010011110010100110111110101111001101110101001 :
(key == 11'b00110101100) ? 46'b1010011101101001000101010101111000100110001101 :
(key == 11'b00110101101) ? 46'b1010011100111101010101010101110111011101110111 :
(key == 11'b00110101110) ? 46'b1010011100010001100111010101110110010101100110 :
(key == 11'b00110101111) ? 46'b1010011011100101111011110101110101001101011011 :
(key == 11'b00110110000) ? 46'b1010011010111010010010010101110100000101010101 :
(key == 11'b00110110001) ? 46'b1010011010001110101011010101110010111101010110 :
(key == 11'b00110110010) ? 46'b1010011001100011000110110101110001110101011100 :
(key == 11'b00110110011) ? 46'b1010011000110111100100010101110000101101100111 :
(key == 11'b00110110100) ? 46'b1010011000001100000011110101101111100101111000 :
(key == 11'b00110110101) ? 46'b1010010111100000100101110101101110011110001110 :
(key == 11'b00110110110) ? 46'b1010010110110101001001110101101101010110101010 :
(key == 11'b00110110111) ? 46'b1010010110001001110000010101101100001111001011 :
(key == 11'b00110111000) ? 46'b1010010101011110011000110101101011000111110010 :
(key == 11'b00110111001) ? 46'b1010010100110011000011110101101010000000011111 :
(key == 11'b00110111010) ? 46'b1010010100000111110000110101101000111001010000 :
(key == 11'b00110111011) ? 46'b1010010011011100100000010101100111110010001000 :
(key == 11'b00110111100) ? 46'b1010010010110001010001110101100110101011000101 :
(key == 11'b00110111101) ? 46'b1010010010000110000101110101100101100100001000 :
(key == 11'b00110111110) ? 46'b1010010001011010111011110101100100011101001111 :
(key == 11'b00110111111) ? 46'b1010010000101111110011110101100011010110011100 :
(key == 11'b00111000000) ? 46'b1010010000000100101110010101100010001111101111 :
(key == 11'b00111000001) ? 46'b1010001111011001101010110101100001001001000111 :
(key == 11'b00111000010) ? 46'b1010001110101110101001110101100000000010100101 :
(key == 11'b00111000011) ? 46'b1010001110000011101010110101011110111100001000 :
(key == 11'b00111000100) ? 46'b1010001101011000101101110101011101110101110000 :
(key == 11'b00111000101) ? 46'b1010001100101101110011010101011100101111011110 :
(key == 11'b00111000110) ? 46'b1010001100000010111010110101011011101001010001 :
(key == 11'b00111000111) ? 46'b1010001011011000000100110101011010100011001010 :
(key == 11'b00111001000) ? 46'b1010001010101101010000110101011001011101001000 :
(key == 11'b00111001001) ? 46'b1010001010000010011110110101011000010111001011 :
(key == 11'b00111001010) ? 46'b1010001001010111101111010101010111010001010100 :
(key == 11'b00111001011) ? 46'b1010001000101101000001110101010110001011100010 :
(key == 11'b00111001100) ? 46'b1010001000000010010110010101010101000101110101 :
(key == 11'b00111001101) ? 46'b1010000111010111101101010101010100000000001110 :
(key == 11'b00111001110) ? 46'b1010000110101101000110010101010010111010101011 :
(key == 11'b00111001111) ? 46'b1010000110000010100001110101010001110101001111 :
(key == 11'b00111010000) ? 46'b1010000101010111111111010101010000101111111000 :
(key == 11'b00111010001) ? 46'b1010000100101101011110110101001111101010100110 :
(key == 11'b00111010010) ? 46'b1010000100000011000000010101001110100101011001 :
(key == 11'b00111010011) ? 46'b1010000011011000100100010101001101100000010001 :
(key == 11'b00111010100) ? 46'b1010000010101110001010010101001100011011001111 :
(key == 11'b00111010101) ? 46'b1010000010000011110010110101001011010110010010 :
(key == 11'b00111010110) ? 46'b1010000001011001011101010101001010010001011011 :
(key == 11'b00111010111) ? 46'b1010000000101111001001110101001001001100101000 :
(key == 11'b00111011000) ? 46'b1010000000000100111000010101001000000111111011 :
(key == 11'b00111011001) ? 46'b1001111111011010101001010101000111000011010011 :
(key == 11'b00111011010) ? 46'b1001111110110000011100010101000101111110110000 :
(key == 11'b00111011011) ? 46'b1001111110000110010001010101000100111010010011 :
(key == 11'b00111011100) ? 46'b1001111101011100001000010101000011110101111010 :
(key == 11'b00111011101) ? 46'b1001111100110010000001110101000010110001100111 :
(key == 11'b00111011110) ? 46'b1001111100000111111101010101000001101101011001 :
(key == 11'b00111011111) ? 46'b1001111011011101111010110101000000101001010000 :
(key == 11'b00111100000) ? 46'b1001111010110011111010110100111111100101001101 :
(key == 11'b00111100001) ? 46'b1001111010001001111100110100111110100001001110 :
(key == 11'b00111100010) ? 46'b1001111001100000000000110100111101011101010101 :
(key == 11'b00111100011) ? 46'b1001111000110110000110110100111100011001100001 :
(key == 11'b00111100100) ? 46'b1001111000001100001111010100111011010101110010 :
(key == 11'b00111100101) ? 46'b1001110111100010011001010100111010010010001000 :
(key == 11'b00111100110) ? 46'b1001110110111000100101110100111001001110100011 :
(key == 11'b00111100111) ? 46'b1001110110001110110100110100111000001011000100 :
(key == 11'b00111101000) ? 46'b1001110101100101000101010100110111000111101001 :
(key == 11'b00111101001) ? 46'b1001110100111011011000010100110110000100010100 :
(key == 11'b00111101010) ? 46'b1001110100010001101100110100110101000001000011 :
(key == 11'b00111101011) ? 46'b1001110011101000000011110100110011111101111000 :
(key == 11'b00111101100) ? 46'b1001110010111110011101010100110010111010110010 :
(key == 11'b00111101101) ? 46'b1001110010010100111000010100110001110111110001 :
(key == 11'b00111101110) ? 46'b1001110001101011010101110100110000110100110101 :
(key == 11'b00111101111) ? 46'b1001110001000001110101010100101111110001111110 :
(key == 11'b00111110000) ? 46'b1001110000011000010110010100101110101111001011 :
(key == 11'b00111110001) ? 46'b1001101111101110111010010100101101101100011111 :
(key == 11'b00111110010) ? 46'b1001101111000101011111110100101100101001110111 :
(key == 11'b00111110011) ? 46'b1001101110011100000111010100101011100111010100 :
(key == 11'b00111110100) ? 46'b1001101101110010110001010100101010100100110110 :
(key == 11'b00111110101) ? 46'b1001101101001001011101010100101001100010011110 :
(key == 11'b00111110110) ? 46'b1001101100100000001011010100101000100000001010 :
(key == 11'b00111110111) ? 46'b1001101011110110111011010100100111011101111011 :
(key == 11'b00111111000) ? 46'b1001101011001101101101010100100110011011110001 :
(key == 11'b00111111001) ? 46'b1001101010100100100001010100100101011001101100 :
(key == 11'b00111111010) ? 46'b1001101001111011010111110100100100010111101100 :
(key == 11'b00111111011) ? 46'b1001101001010010001111110100100011010101110001 :
(key == 11'b00111111100) ? 46'b1001101000101001001010010100100010010011111011 :
(key == 11'b00111111101) ? 46'b1001101000000000000110110100100001010010001010 :
(key == 11'b00111111110) ? 46'b1001100111010111000101010100100000010000011110 :
(key == 11'b00111111111) ? 46'b1001100110101110000101110100011111001110110111 :
(key == 11'b01000000000) ? 46'b1001100110000101001000010100011110001101010100 :
(key == 11'b01000000001) ? 46'b1001100101011100001100110100011101001011110111 :
(key == 11'b01000000010) ? 46'b1001100100110011010011010100011100001010011110 :
(key == 11'b01000000011) ? 46'b1001100100001010011100010100011011001001001011 :
(key == 11'b01000000100) ? 46'b1001100011100001100110110100011010000111111100 :
(key == 11'b01000000101) ? 46'b1001100010111000110011110100011001000110110011 :
(key == 11'b01000000110) ? 46'b1001100010010000000010010100011000000101101101 :
(key == 11'b01000000111) ? 46'b1001100001100111010011010100010111000100101101 :
(key == 11'b01000001000) ? 46'b1001100000111110100110010100010110000011110010 :
(key == 11'b01000001001) ? 46'b1001100000010101111011010100010101000010111100 :
(key == 11'b01000001010) ? 46'b1001011111101101010001110100010100000010001010 :
(key == 11'b01000001011) ? 46'b1001011111000100101010110100010011000001011101 :
(key == 11'b01000001100) ? 46'b1001011110011100000101110100010010000000110101 :
(key == 11'b01000001101) ? 46'b1001011101110011100010110100010001000000010010 :
(key == 11'b01000001110) ? 46'b1001011101001011000001110100001111111111110100 :
(key == 11'b01000001111) ? 46'b1001011100100010100010110100001110111111011011 :
(key == 11'b01000010000) ? 46'b1001011011111010000101110100001101111111000110 :
(key == 11'b01000010001) ? 46'b1001011011010001101010110100001100111110110110 :
(key == 11'b01000010010) ? 46'b1001011010101001010001110100001011111110101011 :
(key == 11'b01000010011) ? 46'b1001011010000000111011010100001010111110100101 :
(key == 11'b01000010100) ? 46'b1001011001011000100110010100001001111110100100 :
(key == 11'b01000010101) ? 46'b1001011000110000010011010100001000111110100111 :
(key == 11'b01000010110) ? 46'b1001011000001000000010010100000111111110101111 :
(key == 11'b01000010111) ? 46'b1001010111011111110011010100000110111110111100 :
(key == 11'b01000011000) ? 46'b1001010110110111100110010100000101111111001101 :
(key == 11'b01000011001) ? 46'b1001010110001111011011010100000100111111100011 :
(key == 11'b01000011010) ? 46'b1001010101100111010010010100000011111111111110 :
(key == 11'b01000011011) ? 46'b1001010100111111001011010100000011000000011110 :
(key == 11'b01000011100) ? 46'b1001010100010111000110010100000010000001000010 :
(key == 11'b01000011101) ? 46'b1001010011101111000011010100000001000001101011 :
(key == 11'b01000011110) ? 46'b1001010011000111000010010100000000000010011001 :
(key == 11'b01000011111) ? 46'b1001010010011111000011010011111111000011001100 :
(key == 11'b01000100000) ? 46'b1001010001110111000101110011111110000100000010 :
(key == 11'b01000100001) ? 46'b1001010001001111001010110011111101000100111110 :
(key == 11'b01000100010) ? 46'b1001010000100111010001110011111100000101111111 :
(key == 11'b01000100011) ? 46'b1001001111111111011010010011111011000111000100 :
(key == 11'b01000100100) ? 46'b1001001111010111100101010011111010001000001110 :
(key == 11'b01000100101) ? 46'b1001001110101111110001110011111001001001011100 :
(key == 11'b01000100110) ? 46'b1001001110001000000000110011111000001010110000 :
(key == 11'b01000100111) ? 46'b1001001101100000010001010011110111001100000111 :
(key == 11'b01000101000) ? 46'b1001001100111000100011110011110110001101100011 :
(key == 11'b01000101001) ? 46'b1001001100010000111000010011110101001111000100 :
(key == 11'b01000101010) ? 46'b1001001011101001001110110011110100010000101010 :
(key == 11'b01000101011) ? 46'b1001001011000001100111010011110011010010010100 :
(key == 11'b01000101100) ? 46'b1001001010011010000001110011110010010100000011 :
(key == 11'b01000101101) ? 46'b1001001001110010011110010011110001010101110110 :
(key == 11'b01000101110) ? 46'b1001001001001010111100010011110000010111101110 :
(key == 11'b01000101111) ? 46'b1001001000100011011100110011101111011001101011 :
(key == 11'b01000110000) ? 46'b1001000111111011111110110011101110011011101011 :
(key == 11'b01000110001) ? 46'b1001000111010100100010110011101101011101110001 :
(key == 11'b01000110010) ? 46'b1001000110101101001000110011101100011111111011 :
(key == 11'b01000110011) ? 46'b1001000110000101110000110011101011100010001010 :
(key == 11'b01000110100) ? 46'b1001000101011110011010110011101010100100011101 :
(key == 11'b01000110101) ? 46'b1001000100110111000110110011101001100110110101 :
(key == 11'b01000110110) ? 46'b1001000100001111110100010011101000101001010001 :
(key == 11'b01000110111) ? 46'b1001000011101000100011110011100111101011110010 :
(key == 11'b01000111000) ? 46'b1001000011000001010101110011100110101110011000 :
(key == 11'b01000111001) ? 46'b1001000010011010001001010011100101110001000001 :
(key == 11'b01000111010) ? 46'b1001000001110010111110110011100100110011110000 :
(key == 11'b01000111011) ? 46'b1001000001001011110101110011100011110110100010 :
(key == 11'b01000111100) ? 46'b1001000000100100101111010011100010111001011010 :
(key == 11'b01000111101) ? 46'b1000111111111101101010010011100001111100010101 :
(key == 11'b01000111110) ? 46'b1000111111010110100111010011100000111111010110 :
(key == 11'b01000111111) ? 46'b1000111110101111100110010011100000000010011010 :
(key == 11'b01001000000) ? 46'b1000111110001000100111010011011111000101100100 :
(key == 11'b01001000001) ? 46'b1000111101100001101001110011011110001000110001 :
(key == 11'b01001000010) ? 46'b1000111100111010101110110011011101001100000011 :
(key == 11'b01001000011) ? 46'b1000111100010011110101010011011100001111011010 :
(key == 11'b01001000100) ? 46'b1000111011101100111101110011011011010010110101 :
(key == 11'b01001000101) ? 46'b1000111011000110001000010011011010010110010100 :
(key == 11'b01001000110) ? 46'b1000111010011111010100010011011001011001111000 :
(key == 11'b01001000111) ? 46'b1000111001111000100010010011011000011101100000 :
(key == 11'b01001001000) ? 46'b1000111001010001110010010011010111100001001100 :
(key == 11'b01001001001) ? 46'b1000111000101011000100010011010110100100111101 :
(key == 11'b01001001010) ? 46'b1000111000000100011000010011010101101000110011 :
(key == 11'b01001001011) ? 46'b1000110111011101101101110011010100101100101101 :
(key == 11'b01001001100) ? 46'b1000110110110111000101010011010011110000101011 :
(key == 11'b01001001101) ? 46'b1000110110010000011110110011010010110100101101 :
(key == 11'b01001001110) ? 46'b1000110101101001111010010011010001111000110100 :
(key == 11'b01001001111) ? 46'b1000110101000011010111010011010000111100111111 :
(key == 11'b01001010000) ? 46'b1000110100011100110110010011010000000001001111 :
(key == 11'b01001010001) ? 46'b1000110011110110010111010011001111000101100011 :
(key == 11'b01001010010) ? 46'b1000110011001111111001110011001110001001111011 :
(key == 11'b01001010011) ? 46'b1000110010101001011110010011001101001110010111 :
(key == 11'b01001010100) ? 46'b1000110010000011000100110011001100010010111000 :
(key == 11'b01001010101) ? 46'b1000110001011100101101010011001011010111011110 :
(key == 11'b01001010110) ? 46'b1000110000110110010111010011001010011100000111 :
(key == 11'b01001010111) ? 46'b1000110000010000000011110011001001100000110101 :
(key == 11'b01001011000) ? 46'b1000101111101001110001010011001000100101100111 :
(key == 11'b01001011001) ? 46'b1000101111000011100001010011000111101010011110 :
(key == 11'b01001011010) ? 46'b1000101110011101010010110011000110101111011000 :
(key == 11'b01001011011) ? 46'b1000101101110111000110010011000101110100010111 :
(key == 11'b01001011100) ? 46'b1000101101010000111011110011000100111001011011 :
(key == 11'b01001011101) ? 46'b1000101100101010110010110011000011111110100010 :
(key == 11'b01001011110) ? 46'b1000101100000100101011110011000011000011101110 :
(key == 11'b01001011111) ? 46'b1000101011011110100110010011000010001000111101 :
(key == 11'b01001100000) ? 46'b1000101010111000100011010011000001001110010010 :
(key == 11'b01001100001) ? 46'b1000101010010010100001110011000000010011101011 :
(key == 11'b01001100010) ? 46'b1000101001101100100001110010111111011001000111 :
(key == 11'b01001100011) ? 46'b1000101001000110100011110010111110011110101000 :
(key == 11'b01001100100) ? 46'b1000101000100000100111110010111101100100001101 :
(key == 11'b01001100101) ? 46'b1000100111111010101101110010111100101001110111 :
(key == 11'b01001100110) ? 46'b1000100111010100110101010010111011101111100100 :
(key == 11'b01001100111) ? 46'b1000100110101110111110110010111010110101010110 :
(key == 11'b01001101000) ? 46'b1000100110001001001001110010111001111011001100 :
(key == 11'b01001101001) ? 46'b1000100101100011010110110010111001000001000110 :
(key == 11'b01001101010) ? 46'b1000100100111101100101110010111000000111000100 :
(key == 11'b01001101011) ? 46'b1000100100010111110110110010110111001101000111 :
(key == 11'b01001101100) ? 46'b1000100011110010001001010010110110010011001110 :
(key == 11'b01001101101) ? 46'b1000100011001100011101010010110101011001011001 :
(key == 11'b01001101110) ? 46'b1000100010100110110011010010110100011111100111 :
(key == 11'b01001101111) ? 46'b1000100010000001001011010010110011100101111011 :
(key == 11'b01001110000) ? 46'b1000100001011011100101010010110010101100010011 :
(key == 11'b01001110001) ? 46'b1000100000110110000000110010110001110010101110 :
(key == 11'b01001110010) ? 46'b1000100000010000011101110010110000111001001101 :
(key == 11'b01001110011) ? 46'b1000011111101010111101010010101111111111110001 :
(key == 11'b01001110100) ? 46'b1000011111000101011101110010101111000110011001 :
(key == 11'b01001110101) ? 46'b1000011110100000000000110010101110001101000101 :
(key == 11'b01001110110) ? 46'b1000011101111010100101010010101101010011110101 :
(key == 11'b01001110111) ? 46'b1000011101010101001011010010101100011010101001 :
(key == 11'b01001111000) ? 46'b1000011100101111110011010010101011100001100001 :
(key == 11'b01001111001) ? 46'b1000011100001010011101010010101010101000011110 :
(key == 11'b01001111010) ? 46'b1000011011100101001000110010101001101111011110 :
(key == 11'b01001111011) ? 46'b1000011010111111110110010010101000110110100010 :
(key == 11'b01001111100) ? 46'b1000011010011010100101110010100111111101101100 :
(key == 11'b01001111101) ? 46'b1000011001110101010110010010100111000100110111 :
(key == 11'b01001111110) ? 46'b1000011001010000001001010010100110001100001001 :
(key == 11'b01001111111) ? 46'b1000011000101010111101110010100101010011011101 :
(key == 11'b01010000000) ? 46'b1000011000000101110011110010100100011010110110 :
(key == 11'b01010000001) ? 46'b1000010111100000101100010010100011100010010011 :
(key == 11'b01010000010) ? 46'b1000010110111011100101110010100010101001110100 :
(key == 11'b01010000011) ? 46'b1000010110010110100001010010100001110001011000 :
(key == 11'b01010000100) ? 46'b1000010101110001011110110010100000111001000010 :
(key == 11'b01010000101) ? 46'b1000010101001100011101110010100000000000101110 :
(key == 11'b01010000110) ? 46'b1000010100100111011110110010011111001000100000 :
(key == 11'b01010000111) ? 46'b1000010100000010100001010010011110010000010100 :
(key == 11'b01010001000) ? 46'b1000010011011101100101110010011101011000001110 :
(key == 11'b01010001001) ? 46'b1000010010111000101011110010011100100000001010 :
(key == 11'b01010001010) ? 46'b1000010010010011110011110010011011101000001011 :
(key == 11'b01010001011) ? 46'b1000010001101110111101010010011010110000010000 :
(key == 11'b01010001100) ? 46'b1000010001001010001000110010011001111000011001 :
(key == 11'b01010001101) ? 46'b1000010000100101010101110010011001000000100110 :
(key == 11'b01010001110) ? 46'b1000010000000000100100110010011000001000110111 :
(key == 11'b01010001111) ? 46'b1000001111011011110101010010010111010001001100 :
(key == 11'b01010010000) ? 46'b1000001110110111000111110010010110011001100101 :
(key == 11'b01010010001) ? 46'b1000001110010010011011110010010101100010000001 :
(key == 11'b01010010010) ? 46'b1000001101101101110001010010010100101010100001 :
(key == 11'b01010010011) ? 46'b1000001101001001001000110010010011110011000110 :
(key == 11'b01010010100) ? 46'b1000001100100100100010010010010010111011101111 :
(key == 11'b01010010101) ? 46'b1000001011111111111101010010010010000100011011 :
(key == 11'b01010010110) ? 46'b1000001011011011011001110010010001001101001011 :
(key == 11'b01010010111) ? 46'b1000001010110110111000010010010000010110000000 :
(key == 11'b01010011000) ? 46'b1000001010010010011000110010001111011110111000 :
(key == 11'b01010011001) ? 46'b1000001001101101111010010010001110100111110100 :
(key == 11'b01010011010) ? 46'b1000001001001001011110010010001101110000110100 :
(key == 11'b01010011011) ? 46'b1000001000100101000011010010001100111001110111 :
(key == 11'b01010011100) ? 46'b1000001000000000101010010010001100000010111111 :
(key == 11'b01010011101) ? 46'b1000000111011100010011010010001011001100001011 :
(key == 11'b01010011110) ? 46'b1000000110110111111101110010001010010101011011 :
(key == 11'b01010011111) ? 46'b1000000110010011101001110010001001011110101110 :
(key == 11'b01010100000) ? 46'b1000000101101111010111110010001000101000000101 :
(key == 11'b01010100001) ? 46'b1000000101001011000111010010000111110001100000 :
(key == 11'b01010100010) ? 46'b1000000100100110111000110010000110111010111111 :
(key == 11'b01010100011) ? 46'b1000000100000010101011110010000110000100100010 :
(key == 11'b01010100100) ? 46'b1000000011011110100000010010000101001110001000 :
(key == 11'b01010100101) ? 46'b1000000010111010010110110010000100010111110010 :
(key == 11'b01010100110) ? 46'b1000000010010110001110110010000011100001100001 :
(key == 11'b01010100111) ? 46'b1000000001110010001000110010000010101011010011 :
(key == 11'b01010101000) ? 46'b1000000001001110000100010010000001110101001001 :
(key == 11'b01010101001) ? 46'b1000000000101010000001010010000000111111000010 :
(key == 11'b01010101010) ? 46'b1000000000000110000000010010000000001001000000 :
(key == 11'b01010101011) ? 46'b0111111111100010000000110001111111010011000001 :
(key == 11'b01010101100) ? 46'b0111111110111110000011010001111110011101000110 :
(key == 11'b01010101101) ? 46'b0111111110011010000111010001111101100111001111 :
(key == 11'b01010101110) ? 46'b0111111101110110001100110001111100110001011100 :
(key == 11'b01010101111) ? 46'b0111111101010010010011110001111011111011101100 :
(key == 11'b01010110000) ? 46'b0111111100101110011100110001111011000110000000 :
(key == 11'b01010110001) ? 46'b0111111100001010100111110001111010010000011000 :
(key == 11'b01010110010) ? 46'b0111111011100110110011110001111001011010110100 :
(key == 11'b01010110011) ? 46'b0111111011000011000001110001111000100101010011 :
(key == 11'b01010110100) ? 46'b0111111010011111010001110001110111101111110111 :
(key == 11'b01010110101) ? 46'b0111111001111011100010110001110110111010011101 :
(key == 11'b01010110110) ? 46'b0111111001010111110101110001110110000101001000 :
(key == 11'b01010110111) ? 46'b0111111000110100001010110001110101001111110111 :
(key == 11'b01010111000) ? 46'b0111111000010000100000110001110100011010101000 :
(key == 11'b01010111001) ? 46'b0111110111101100111000110001110011100101011110 :
(key == 11'b01010111010) ? 46'b0111110111001001010010110001110010110000011000 :
(key == 11'b01010111011) ? 46'b0111110110100101101101110001110001111011010101 :
(key == 11'b01010111100) ? 46'b0111110110000010001010110001110001000110010110 :
(key == 11'b01010111101) ? 46'b0111110101011110101001010001110000010001011011 :
(key == 11'b01010111110) ? 46'b0111110100111011001001110001101111011100100011 :
(key == 11'b01010111111) ? 46'b0111110100010111101011110001101110100111110000 :
(key == 11'b01011000000) ? 46'b0111110011110100001111010001101101110010111111 :
(key == 11'b01011000001) ? 46'b0111110011010000110100110001101100111110010011 :
(key == 11'b01011000010) ? 46'b0111110010101101011011010001101100001001101010 :
(key == 11'b01011000011) ? 46'b0111110010001010000011110001101011010101000100 :
(key == 11'b01011000100) ? 46'b0111110001100110101110010001101010100000100011 :
(key == 11'b01011000101) ? 46'b0111110001000011011001110001101001101100000101 :
(key == 11'b01011000110) ? 46'b0111110000100000000111010001101000110111101011 :
(key == 11'b01011000111) ? 46'b0111101111111100110110010001101000000011010100 :
(key == 11'b01011001000) ? 46'b0111101111011001100111010001100111001111000001 :
(key == 11'b01011001001) ? 46'b0111101110110110011001010001100110011010110010 :
(key == 11'b01011001010) ? 46'b0111101110010011001101010001100101100110100110 :
(key == 11'b01011001011) ? 46'b0111101101110000000011010001100100110010011110 :
(key == 11'b01011001100) ? 46'b0111101101001100111010010001100011111110011010 :
(key == 11'b01011001101) ? 46'b0111101100101001110011010001100011001010011001 :
(key == 11'b01011001110) ? 46'b0111101100000110101101110001100010010110011100 :
(key == 11'b01011001111) ? 46'b0111101011100011101001110001100001100010100010 :
(key == 11'b01011010000) ? 46'b0111101011000000100111010001100000101110101011 :
(key == 11'b01011010001) ? 46'b0111101010011101100110110001011111111010111001 :
(key == 11'b01011010010) ? 46'b0111101001111010100111110001011111000111001010 :
(key == 11'b01011010011) ? 46'b0111101001010111101010010001011110010011011111 :
(key == 11'b01011010100) ? 46'b0111101000110100101110110001011101011111111000 :
(key == 11'b01011010101) ? 46'b0111101000010001110100010001011100101100010011 :
(key == 11'b01011010110) ? 46'b0111100111101110111011110001011011111000110011 :
(key == 11'b01011010111) ? 46'b0111100111001100000100110001011011000101010110 :
(key == 11'b01011011000) ? 46'b0111100110101001001111010001011010010001111100 :
(key == 11'b01011011001) ? 46'b0111100110000110011011110001011001011110100111 :
(key == 11'b01011011010) ? 46'b0111100101100011101001110001011000101011010100 :
(key == 11'b01011011011) ? 46'b0111100101000000111000110001010111111000000101 :
(key == 11'b01011011100) ? 46'b0111100100011110001010010001010111000100111010 :
(key == 11'b01011011101) ? 46'b0111100011111011011100110001010110010001110010 :
(key == 11'b01011011110) ? 46'b0111100011011000110000110001010101011110101110 :
(key == 11'b01011011111) ? 46'b0111100010110110000110110001010100101011101101 :
(key == 11'b01011100000) ? 46'b0111100010010011011110010001010011111000110000 :
(key == 11'b01011100001) ? 46'b0111100001110000110111010001010011000101110111 :
(key == 11'b01011100010) ? 46'b0111100001001110010001110001010010010011000000 :
(key == 11'b01011100011) ? 46'b0111100000101011101110010001010001100000001110 :
(key == 11'b01011100100) ? 46'b0111100000001001001011110001010000101101011111 :
(key == 11'b01011100101) ? 46'b0111011111100110101011010001001111111010110011 :
(key == 11'b01011100110) ? 46'b0111011111000100001100010001001111001000001011 :
(key == 11'b01011100111) ? 46'b0111011110100001101110110001001110010101100110 :
(key == 11'b01011101000) ? 46'b0111011101111111010010110001001101100011000101 :
(key == 11'b01011101001) ? 46'b0111011101011100111000010001001100110000100111 :
(key == 11'b01011101010) ? 46'b0111011100111010011111110001001011111110001101 :
(key == 11'b01011101011) ? 46'b0111011100011000001000110001001011001011110110 :
(key == 11'b01011101100) ? 46'b0111011011110101110010110001001010011001100011 :
(key == 11'b01011101101) ? 46'b0111011011010011011110110001001001100111010011 :
(key == 11'b01011101110) ? 46'b0111011010110001001100110001001000110101000111 :
(key == 11'b01011101111) ? 46'b0111011010001110111011110001001000000010111110 :
(key == 11'b01011110000) ? 46'b0111011001101100101100010001000111010000111000 :
(key == 11'b01011110001) ? 46'b0111011001001010011110110001000110011110110110 :
(key == 11'b01011110010) ? 46'b0111011000101000010010010001000101101100110111 :
(key == 11'b01011110011) ? 46'b0111011000000110000111110001000100111010111100 :
(key == 11'b01011110100) ? 46'b0111010111100011111110110001000100001001000100 :
(key == 11'b01011110101) ? 46'b0111010111000001110111010001000011010111001111 :
(key == 11'b01011110110) ? 46'b0111010110011111110001010001000010100101011110 :
(key == 11'b01011110111) ? 46'b0111010101111101101100110001000001110011110001 :
(key == 11'b01011111000) ? 46'b0111010101011011101010010001000001000010000111 :
(key == 11'b01011111001) ? 46'b0111010100111001101000110001000000010000100000 :
(key == 11'b01011111010) ? 46'b0111010100010111101001010000111111011110111101 :
(key == 11'b01011111011) ? 46'b0111010011110101101010110000111110101101011100 :
(key == 11'b01011111100) ? 46'b0111010011010011101110010000111101111011111111 :
(key == 11'b01011111101) ? 46'b0111010010110001110011010000111101001010100110 :
(key == 11'b01011111110) ? 46'b0111010010001111111001110000111100011001010000 :
(key == 11'b01011111111) ? 46'b0111010001101110000001110000111011100111111110 :
(key == 11'b01100000000) ? 46'b0111010001001100001011010000111010110110101111 :
(key == 11'b01100000001) ? 46'b0111010000101010010110010000111010000101100011 :
(key == 11'b01100000010) ? 46'b0111010000001000100010110000111001010100011010 :
(key == 11'b01100000011) ? 46'b0111001111100110110000110000111000100011010101 :
(key == 11'b01100000100) ? 46'b0111001111000101000000010000110111110010010010 :
(key == 11'b01100000101) ? 46'b0111001110100011010001110000110111000001010100 :
(key == 11'b01100000110) ? 46'b0111001110000001100100010000110110010000011001 :
(key == 11'b01100000111) ? 46'b0111001101011111111000110000110101011111100001 :
(key == 11'b01100001000) ? 46'b0111001100111110001110010000110100101110101100 :
(key == 11'b01100001001) ? 46'b0111001100011100100101110000110011111101111011 :
(key == 11'b01100001010) ? 46'b0111001011111010111110110000110011001101001110 :
(key == 11'b01100001011) ? 46'b0111001011011001011000110000110010011100100011 :
(key == 11'b01100001100) ? 46'b0111001010110111110100110000110001101011111100 :
(key == 11'b01100001101) ? 46'b0111001010010110010010010000110000111011011000 :
(key == 11'b01100001110) ? 46'b0111001001110100110001010000110000001010110111 :
(key == 11'b01100001111) ? 46'b0111001001010011010001010000101111011010011001 :
(key == 11'b01100010000) ? 46'b0111001000110001110011010000101110101001111111 :
(key == 11'b01100010001) ? 46'b0111001000010000010110110000101101111001101000 :
(key == 11'b01100010010) ? 46'b0111000111101110111011110000101101001001010101 :
(key == 11'b01100010011) ? 46'b0111000111001101100010010000101100011001000101 :
(key == 11'b01100010100) ? 46'b0111000110101100001010010000101011101000111000 :
(key == 11'b01100010101) ? 46'b0111000110001010110011110000101010111000101110 :
(key == 11'b01100010110) ? 46'b0111000101101001011110110000101010001000100111 :
(key == 11'b01100010111) ? 46'b0111000101001000001011010000101001011000100100 :
(key == 11'b01100011000) ? 46'b0111000100100110111001010000101000101000100100 :
(key == 11'b01100011001) ? 46'b0111000100000101101000110000100111111000100111 :
(key == 11'b01100011010) ? 46'b0111000011100100011001110000100111001000101110 :
(key == 11'b01100011011) ? 46'b0111000011000011001100010000100110011000111000 :
(key == 11'b01100011100) ? 46'b0111000010100010000000010000100101101001000101 :
(key == 11'b01100011101) ? 46'b0111000010000000110101110000100100111001010101 :
(key == 11'b01100011110) ? 46'b0111000001011111101100010000100100001001100111 :
(key == 11'b01100011111) ? 46'b0111000000111110100100110000100011011001111110 :
(key == 11'b01100100000) ? 46'b0111000000011101011110110000100010101010011000 :
(key == 11'b01100100001) ? 46'b0110111111111100011010010000100001111010110101 :
(key == 11'b01100100010) ? 46'b0110111111011011010111010000100001001011010101 :
(key == 11'b01100100011) ? 46'b0110111110111010010101110000100000011011111001 :
(key == 11'b01100100100) ? 46'b0110111110011001010101010000011111101100011111 :
(key == 11'b01100100101) ? 46'b0110111101111000010110110000011110111101001001 :
(key == 11'b01100100110) ? 46'b0110111101010111011001110000011110001101110110 :
(key == 11'b01100100111) ? 46'b0110111100110110011101110000011101011110100110 :
(key == 11'b01100101000) ? 46'b0110111100010101100011110000011100101111011010 :
(key == 11'b01100101001) ? 46'b0110111011110100101010110000011100000000010000 :
(key == 11'b01100101010) ? 46'b0110111011010011110011110000011011010001001010 :
(key == 11'b01100101011) ? 46'b0110111010110010111101110000011010100010000110 :
(key == 11'b01100101100) ? 46'b0110111010010010001001110000011001110011000111 :
(key == 11'b01100101101) ? 46'b0110111001110001010110110000011001000100001010 :
(key == 11'b01100101110) ? 46'b0110111001010000100101010000011000010101010000 :
(key == 11'b01100101111) ? 46'b0110111000101111110101010000010111100110011001 :
(key == 11'b01100110000) ? 46'b0110111000001111000110110000010110110111100110 :
(key == 11'b01100110001) ? 46'b0110110111101110011001110000010110001000110101 :
(key == 11'b01100110010) ? 46'b0110110111001101101110010000010101011010001000 :
(key == 11'b01100110011) ? 46'b0110110110101101000100010000010100101011011110 :
(key == 11'b01100110100) ? 46'b0110110110001100011011110000010011111100111000 :
(key == 11'b01100110101) ? 46'b0110110101101011110100010000010011001110010011 :
(key == 11'b01100110110) ? 46'b0110110101001011001110110000010010011111110011 :
(key == 11'b01100110111) ? 46'b0110110100101010101010010000010001110001010101 :
(key == 11'b01100111000) ? 46'b0110110100001010000111110000010001000010111011 :
(key == 11'b01100111001) ? 46'b0110110011101001100110010000010000010100100011 :
(key == 11'b01100111010) ? 46'b0110110011001001000110010000001111100110001111 :
(key == 11'b01100111011) ? 46'b0110110010101000100111110000001110110111111110 :
(key == 11'b01100111100) ? 46'b0110110010001000001010110000001110001001110000 :
(key == 11'b01100111101) ? 46'b0110110001100111101111010000001101011011100101 :
(key == 11'b01100111110) ? 46'b0110110001000111010101010000001100101101011101 :
(key == 11'b01100111111) ? 46'b0110110000100110111100010000001011111111011000 :
(key == 11'b01101000000) ? 46'b0110110000000110100101010000001011010001010110 :
(key == 11'b01101000001) ? 46'b0110101111100110001111010000001010100011010111 :
(key == 11'b01101000010) ? 46'b0110101111000101111010110000001001110101011100 :
(key == 11'b01101000011) ? 46'b0110101110100101100111110000001001000111100011 :
(key == 11'b01101000100) ? 46'b0110101110000101010110010000001000011001101101 :
(key == 11'b01101000101) ? 46'b0110101101100101000110010000000111101011111011 :
(key == 11'b01101000110) ? 46'b0110101101000100110111110000000110111110001100 :
(key == 11'b01101000111) ? 46'b0110101100100100101010010000000110010000011111 :
(key == 11'b01101001000) ? 46'b0110101100000100011110110000000101100010110110 :
(key == 11'b01101001001) ? 46'b0110101011100100010100010000000100110101001111 :
(key == 11'b01101001010) ? 46'b0110101011000100001011010000000100000111101100 :
(key == 11'b01101001011) ? 46'b0110101010100100000011110000000011011010001100 :
(key == 11'b01101001100) ? 46'b0110101010000011111101110000000010101100101111 :
(key == 11'b01101001101) ? 46'b0110101001100011111001010000000001111111010101 :
(key == 11'b01101001110) ? 46'b0110101001000011110101110000000001010001111101 :
(key == 11'b01101001111) ? 46'b0110101000100011110011110000000000100100101001 :
(key == 11'b01101010000) ? 46'b0110101000000011110011001111111111110111010111 :
(key == 11'b01101010001) ? 46'b0110100111100011110100001111111111001010001001 :
(key == 11'b01101010010) ? 46'b0110100111000011110110101111111110011100111110 :
(key == 11'b01101010011) ? 46'b0110100110100011111010101111111101101111110110 :
(key == 11'b01101010100) ? 46'b0110100110000011111111101111111101000010110000 :
(key == 11'b01101010101) ? 46'b0110100101100100000110001111111100010101101110 :
(key == 11'b01101010110) ? 46'b0110100101000100001110001111111011101000101111 :
(key == 11'b01101010111) ? 46'b0110100100100100010111101111111010111011110010 :
(key == 11'b01101011000) ? 46'b0110100100000100100010101111111010001110111001 :
(key == 11'b01101011001) ? 46'b0110100011100100101110101111111001100010000011 :
(key == 11'b01101011010) ? 46'b0110100011000100111100101111111000110101010000 :
(key == 11'b01101011011) ? 46'b0110100010100101001011101111111000001000011111 :
(key == 11'b01101011100) ? 46'b0110100010000101011100001111110111011011110010 :
(key == 11'b01101011101) ? 46'b0110100001100101101101101111110110101111000111 :
(key == 11'b01101011110) ? 46'b0110100001000110000001001111110110000010011111 :
(key == 11'b01101011111) ? 46'b0110100000100110010101101111110101010101111011 :
(key == 11'b01101100000) ? 46'b0110100000000110101011101111110100101001011001 :
(key == 11'b01101100001) ? 46'b0110011111100111000011001111110011111100111010 :
(key == 11'b01101100010) ? 46'b0110011111000111011011101111110011010000011110 :
(key == 11'b01101100011) ? 46'b0110011110100111110110001111110010100100000101 :
(key == 11'b01101100100) ? 46'b0110011110001000010001101111110001110111101111 :
(key == 11'b01101100101) ? 46'b0110011101101000101110101111110001001011011100 :
(key == 11'b01101100110) ? 46'b0110011101001001001101001111110000011111001100 :
(key == 11'b01101100111) ? 46'b0110011100101001101100101111101111110010111111 :
(key == 11'b01101101000) ? 46'b0110011100001010001101101111101111000110110100 :
(key == 11'b01101101001) ? 46'b0110011011101010110000001111101110011010101101 :
(key == 11'b01101101010) ? 46'b0110011011001011010100001111101101101110101000 :
(key == 11'b01101101011) ? 46'b0110011010101011111001001111101101000010100110 :
(key == 11'b01101101100) ? 46'b0110011010001100011111101111101100010110100111 :
(key == 11'b01101101101) ? 46'b0110011001101101000111101111101011101010101011 :
(key == 11'b01101101110) ? 46'b0110011001001101110001001111101010111110110011 :
(key == 11'b01101101111) ? 46'b0110011000101110011100001111101010010010111101 :
(key == 11'b01101110000) ? 46'b0110011000001111001000001111101001100111001001 :
(key == 11'b01101110001) ? 46'b0110010111101111110101101111101000111011011001 :
(key == 11'b01101110010) ? 46'b0110010111010000100100001111101000001111101011 :
(key == 11'b01101110011) ? 46'b0110010110110001010100101111100111100100000001 :
(key == 11'b01101110100) ? 46'b0110010110010010000110001111100110111000011001 :
(key == 11'b01101110101) ? 46'b0110010101110010111001001111100110001100110100 :
(key == 11'b01101110110) ? 46'b0110010101010011101101001111100101100001010010 :
(key == 11'b01101110111) ? 46'b0110010100110100100011001111100100110101110011 :
(key == 11'b01101111000) ? 46'b0110010100010101011010001111100100001010010110 :
(key == 11'b01101111001) ? 46'b0110010011110110010010001111100011011110111100 :
(key == 11'b01101111010) ? 46'b0110010011010111001100001111100010110011100110 :
(key == 11'b01101111011) ? 46'b0110010010111000000111001111100010001000010010 :
(key == 11'b01101111100) ? 46'b0110010010011001000011101111100001011101000001 :
(key == 11'b01101111101) ? 46'b0110010001111010000001001111100000110001110010 :
(key == 11'b01101111110) ? 46'b0110010001011011000000001111100000000110100111 :
(key == 11'b01101111111) ? 46'b0110010000111100000000101111011111011011011110 :
(key == 11'b01110000000) ? 46'b0110010000011101000010101111011110110000011001 :
(key == 11'b01110000001) ? 46'b0110001111111110000101101111011110000101010101 :
(key == 11'b01110000010) ? 46'b0110001111011111001010001111011101011010010101 :
(key == 11'b01110000011) ? 46'b0110001111000000010000001111011100101111011000 :
(key == 11'b01110000100) ? 46'b0110001110100001010111001111011100000100011101 :
(key == 11'b01110000101) ? 46'b0110001110000010011111101111011011011001100101 :
(key == 11'b01110000110) ? 46'b0110001101100011101001101111011010101110110000 :
(key == 11'b01110000111) ? 46'b0110001101000100110101001111011010000011111110 :
(key == 11'b01110001000) ? 46'b0110001100100110000001101111011001011001001111 :
(key == 11'b01110001001) ? 46'b0110001100000111001111001111011000101110100010 :
(key == 11'b01110001010) ? 46'b0110001011101000011110101111011000000011111000 :
(key == 11'b01110001011) ? 46'b0110001011001001101111001111010111011001010001 :
(key == 11'b01110001100) ? 46'b0110001010101011000001001111010110101110101101 :
(key == 11'b01110001101) ? 46'b0110001010001100010100001111010110000100001011 :
(key == 11'b01110001110) ? 46'b0110001001101101101000101111010101011001101100 :
(key == 11'b01110001111) ? 46'b0110001001001110111110101111010100101111010000 :
(key == 11'b01110010000) ? 46'b0110001000110000010101101111010100000100110110 :
(key == 11'b01110010001) ? 46'b0110001000010001101110001111010011011010100000 :
(key == 11'b01110010010) ? 46'b0110000111110011001000001111010010110000001100 :
(key == 11'b01110010011) ? 46'b0110000111010100100011001111010010000101111011 :
(key == 11'b01110010100) ? 46'b0110000110110101111111101111010001011011101101 :
(key == 11'b01110010101) ? 46'b0110000110010111011101101111010000110001100001 :
(key == 11'b01110010110) ? 46'b0110000101111000111100101111010000000111011000 :
(key == 11'b01110010111) ? 46'b0110000101011010011101001111001111011101010010 :
(key == 11'b01110011000) ? 46'b0110000100111011111110101111001110110011001110 :
(key == 11'b01110011001) ? 46'b0110000100011101100001101111001110001001001101 :
(key == 11'b01110011010) ? 46'b0110000011111111000110001111001101011111010000 :
(key == 11'b01110011011) ? 46'b0110000011100000101100001111001100110101010101 :
(key == 11'b01110011100) ? 46'b0110000011000010010011001111001100001011011100 :
(key == 11'b01110011101) ? 46'b0110000010100011111011001111001011100001100110 :
(key == 11'b01110011110) ? 46'b0110000010000101100100101111001010110111110011 :
(key == 11'b01110011111) ? 46'b0110000001100111001111101111001010001110000010 :
(key == 11'b01110100000) ? 46'b0110000001001000111100001111001001100100010101 :
(key == 11'b01110100001) ? 46'b0110000000101010101001101111001000111010101010 :
(key == 11'b01110100010) ? 46'b0110000000001100011000001111001000010001000001 :
(key == 11'b01110100011) ? 46'b0101111111101110001000001111000111100111011011 :
(key == 11'b01110100100) ? 46'b0101111111001111111001101111000110111101111000 :
(key == 11'b01110100101) ? 46'b0101111110110001101100101111000110010100011000 :
(key == 11'b01110100110) ? 46'b0101111110010011100000101111000101101010111010 :
(key == 11'b01110100111) ? 46'b0101111101110101010101101111000101000001011111 :
(key == 11'b01110101000) ? 46'b0101111101010111001100101111000100011000000111 :
(key == 11'b01110101001) ? 46'b0101111100111001000100001111000011101110110000 :
(key == 11'b01110101010) ? 46'b0101111100011010111101101111000011000101011110 :
(key == 11'b01110101011) ? 46'b0101111011111100111000001111000010011100001101 :
(key == 11'b01110101100) ? 46'b0101111011011110110011101111000001110010111111 :
(key == 11'b01110101101) ? 46'b0101111011000000110000101111000001001001110100 :
(key == 11'b01110101110) ? 46'b0101111010100010101111001111000000100000101100 :
(key == 11'b01110101111) ? 46'b0101111010000100101110101110111111110111100110 :
(key == 11'b01110110000) ? 46'b0101111001100110101111101110111111001110100011 :
(key == 11'b01110110001) ? 46'b0101111001001000110001101110111110100101100010 :
(key == 11'b01110110010) ? 46'b0101111000101010110101001110111101111100100100 :
(key == 11'b01110110011) ? 46'b0101111000001100111010001110111101010011101001 :
(key == 11'b01110110100) ? 46'b0101110111101111000000001110111100101010110000 :
(key == 11'b01110110101) ? 46'b0101110111010001000111001110111100000001111010 :
(key == 11'b01110110110) ? 46'b0101110110110011010000001110111011011001000111 :
(key == 11'b01110110111) ? 46'b0101110110010101011001101110111010110000010110 :
(key == 11'b01110111000) ? 46'b0101110101110111100101001110111010000111101000 :
(key == 11'b01110111001) ? 46'b0101110101011001110001001110111001011110111100 :
(key == 11'b01110111010) ? 46'b0101110100111011111111001110111000110110010011 :
(key == 11'b01110111011) ? 46'b0101110100011110001110001110111000001101101101 :
(key == 11'b01110111100) ? 46'b0101110100000000011110001110110111100101001001 :
(key == 11'b01110111101) ? 46'b0101110011100010101111101110110110111100100111 :
(key == 11'b01110111110) ? 46'b0101110011000101000010001110110110010100001000 :
(key == 11'b01110111111) ? 46'b0101110010100111010110001110110101101011101100 :
(key == 11'b01111000000) ? 46'b0101110010001001101011101110110101000011010011 :
(key == 11'b01111000001) ? 46'b0101110001101100000010001110110100011010111100 :
(key == 11'b01111000010) ? 46'b0101110001001110011010001110110011110010101000 :
(key == 11'b01111000011) ? 46'b0101110000110000110011001110110011001010010110 :
(key == 11'b01111000100) ? 46'b0101110000010011001101001110110010100010000110 :
(key == 11'b01111000101) ? 46'b0101101111110101101000101110110001111001111010 :
(key == 11'b01111000110) ? 46'b0101101111011000000101101110110001010001110000 :
(key == 11'b01111000111) ? 46'b0101101110111010100011101110110000101001101000 :
(key == 11'b01111001000) ? 46'b0101101110011101000011001110110000000001100011 :
(key == 11'b01111001001) ? 46'b0101101101111111100011101110101111011001100001 :
(key == 11'b01111001010) ? 46'b0101101101100010000101101110101110110001100001 :
(key == 11'b01111001011) ? 46'b0101101101000100101000101110101110001001100100 :
(key == 11'b01111001100) ? 46'b0101101100100111001100101110101101100001101001 :
(key == 11'b01111001101) ? 46'b0101101100001001110010101110101100111001110001 :
(key == 11'b01111001110) ? 46'b0101101011101100011001001110101100010001111011 :
(key == 11'b01111001111) ? 46'b0101101011001111000001001110101011101010000111 :
(key == 11'b01111010000) ? 46'b0101101010110001101010101110101011000010010111 :
(key == 11'b01111010001) ? 46'b0101101010010100010101001110101010011010101001 :
(key == 11'b01111010010) ? 46'b0101101001110111000001001110101001110010111101 :
(key == 11'b01111010011) ? 46'b0101101001011001101110001110101001001011010100 :
(key == 11'b01111010100) ? 46'b0101101000111100011100001110101000100011101101 :
(key == 11'b01111010101) ? 46'b0101101000011111001011101110100111111100001001 :
(key == 11'b01111010110) ? 46'b0101101000000001111100101110100111010100101000 :
(key == 11'b01111010111) ? 46'b0101100111100100101110101110100110101101001001 :
(key == 11'b01111011000) ? 46'b0101100111000111100001101110100110000101101100 :
(key == 11'b01111011001) ? 46'b0101100110101010010110001110100101011110010010 :
(key == 11'b01111011010) ? 46'b0101100110001101001011101110100100110110111010 :
(key == 11'b01111011011) ? 46'b0101100101110000000010101110100100001111100101 :
(key == 11'b01111011100) ? 46'b0101100101010010111010101110100011101000010010 :
(key == 11'b01111011101) ? 46'b0101100100110101110100001110100011000001000010 :
(key == 11'b01111011110) ? 46'b0101100100011000101110101110100010011001110101 :
(key == 11'b01111011111) ? 46'b0101100011111011101010101110100001110010101010 :
(key == 11'b01111100000) ? 46'b0101100011011110100111101110100001001011100001 :
(key == 11'b01111100001) ? 46'b0101100011000001100101101110100000100100011010 :
(key == 11'b01111100010) ? 46'b0101100010100100100101001110011111111101010111 :
(key == 11'b01111100011) ? 46'b0101100010000111100110001110011111010110010110 :
(key == 11'b01111100100) ? 46'b0101100001101010101000001110011110101111010111 :
(key == 11'b01111100101) ? 46'b0101100001001101101011001110011110001000011010 :
(key == 11'b01111100110) ? 46'b0101100000110000101111001110011101100001100000 :
(key == 11'b01111100111) ? 46'b0101100000010011110101001110011100111010101001 :
(key == 11'b01111101000) ? 46'b0101011111110110111011101110011100010011110100 :
(key == 11'b01111101001) ? 46'b0101011111011010000011101110011011101101000001 :
(key == 11'b01111101010) ? 46'b0101011110111101001100101110011011000110010001 :
(key == 11'b01111101011) ? 46'b0101011110100000010111001110011010011111100011 :
(key == 11'b01111101100) ? 46'b0101011110000011100011001110011001111000111000 :
(key == 11'b01111101101) ? 46'b0101011101100110101111101110011001010010001111 :
(key == 11'b01111101110) ? 46'b0101011101001001111101101110011000101011101000 :
(key == 11'b01111101111) ? 46'b0101011100101101001101001110011000000101000101 :
(key == 11'b01111110000) ? 46'b0101011100010000011101101110010111011110100011 :
(key == 11'b01111110001) ? 46'b0101011011110011101111001110010110111000000100 :
(key == 11'b01111110010) ? 46'b0101011011010111000010001110010110010001100111 :
(key == 11'b01111110011) ? 46'b0101011010111010010110001110010101101011001101 :
(key == 11'b01111110100) ? 46'b0101011010011101101011001110010101000100110101 :
(key == 11'b01111110101) ? 46'b0101011010000001000001101110010100011110011111 :
(key == 11'b01111110110) ? 46'b0101011001100100011001001110010011111000001100 :
(key == 11'b01111110111) ? 46'b0101011001000111110010001110010011010001111011 :
(key == 11'b01111111000) ? 46'b0101011000101011001100001110010010101011101101 :
(key == 11'b01111111001) ? 46'b0101011000001110100111101110010010000101100001 :
(key == 11'b01111111010) ? 46'b0101010111110010000011101110010001011111010111 :
(key == 11'b01111111011) ? 46'b0101010111010101100001101110010000111001010001 :
(key == 11'b01111111100) ? 46'b0101010110111001000000001110010000010011001100 :
(key == 11'b01111111101) ? 46'b0101010110011100100000001110001111101101001001 :
(key == 11'b01111111110) ? 46'b0101010110000000000001101110001111000111001010 :
(key == 11'b01111111111) ? 46'b0101010101100011100011101110001110100001001100 :
(key == 11'b10000000000) ? 46'b0101010101000111000111101110001101111011010001 :
(key == 11'b10000000001) ? 46'b0101010100101010101100001110001101010101011000 :
(key == 11'b10000000010) ? 46'b0101010100001110010010001110001100101111100001 :
(key == 11'b10000000011) ? 46'b0101010011110001111001001110001100001001101101 :
(key == 11'b10000000100) ? 46'b0101010011010101100001101110001011100011111011 :
(key == 11'b10000000101) ? 46'b0101010010111001001011001110001010111110001100 :
(key == 11'b10000000110) ? 46'b0101010010011100110101101110001010011000011111 :
(key == 11'b10000000111) ? 46'b0101010010000000100001101110001001110010110100 :
(key == 11'b10000001000) ? 46'b0101010001100100001110101110001001001101001100 :
(key == 11'b10000001001) ? 46'b0101010001000111111100101110001000100111100110 :
(key == 11'b10000001010) ? 46'b0101010000101011101100001110001000000010000010 :
(key == 11'b10000001011) ? 46'b0101010000001111011100101110000111011100100001 :
(key == 11'b10000001100) ? 46'b0101001111110011001110001110000110110111000001 :
(key == 11'b10000001101) ? 46'b0101001111010111000001001110000110010001100101 :
(key == 11'b10000001110) ? 46'b0101001110111010110101001110000101101100001010 :
(key == 11'b10000001111) ? 46'b0101001110011110101010001110000101000110110010 :
(key == 11'b10000010000) ? 46'b0101001110000010100000101110000100100001011100 :
(key == 11'b10000010001) ? 46'b0101001101100110011000001110000011111100001001 :
(key == 11'b10000010010) ? 46'b0101001101001010010000101110000011010110111000 :
(key == 11'b10000010011) ? 46'b0101001100101110001010101110000010110001101001 :
(key == 11'b10000010100) ? 46'b0101001100010010000101101110000010001100011101 :
(key == 11'b10000010101) ? 46'b0101001011110110000010001110000001100111010011 :
(key == 11'b10000010110) ? 46'b0101001011011001111111001110000001000010001011 :
(key == 11'b10000010111) ? 46'b0101001010111101111101101110000000011101000101 :
(key == 11'b10000011000) ? 46'b0101001010100001111101101101111111111000000010 :
(key == 11'b10000011001) ? 46'b0101001010000101111110001101111111010011000001 :
(key == 11'b10000011010) ? 46'b0101001001101010000000001101111110101110000010 :
(key == 11'b10000011011) ? 46'b0101001001001110000011101101111110001001000110 :
(key == 11'b10000011100) ? 46'b0101001000110010000111101101111101100100001100 :
(key == 11'b10000011101) ? 46'b0101001000010110001101001101111100111111010100 :
(key == 11'b10000011110) ? 46'b0101000111111010010011101101111100011010011110 :
(key == 11'b10000011111) ? 46'b0101000111011110011011101101111011110101101011 :
(key == 11'b10000100000) ? 46'b0101000111000010100100101101111011010000111011 :
(key == 11'b10000100001) ? 46'b0101000110100110101110101101111010101100001100 :
(key == 11'b10000100010) ? 46'b0101000110001010111001101101111010000111011111 :
(key == 11'b10000100011) ? 46'b0101000101101111000110001101111001100010110101 :
(key == 11'b10000100100) ? 46'b0101000101010011010011101101111000111110001101 :
(key == 11'b10000100101) ? 46'b0101000100110111100010001101111000011001101000 :
(key == 11'b10000100110) ? 46'b0101000100011011110001101101110111110101000100 :
(key == 11'b10000100111) ? 46'b0101000100000000000010101101110111010000100011 :
(key == 11'b10000101000) ? 46'b0101000011100100010100101101110110101100000100 :
(key == 11'b10000101001) ? 46'b0101000011001000101000001101110110000111101000 :
(key == 11'b10000101010) ? 46'b0101000010101100111100001101110101100011001101 :
(key == 11'b10000101011) ? 46'b0101000010010001010001101101110100111110110101 :
(key == 11'b10000101100) ? 46'b0101000001110101101000101101110100011010100000 :
(key == 11'b10000101101) ? 46'b0101000001011010000000001101110011110110001100 :
(key == 11'b10000101110) ? 46'b0101000000111110011001001101110011010001111010 :
(key == 11'b10000101111) ? 46'b0101000000100010110011001101110010101101101011 :
(key == 11'b10000110000) ? 46'b0101000000000111001110001101110010001001011110 :
(key == 11'b10000110001) ? 46'b0100111111101011101010101101110001100101010100 :
(key == 11'b10000110010) ? 46'b0100111111010000000111101101110001000001001011 :
(key == 11'b10000110011) ? 46'b0100111110110100100110001101110000011101000100 :
(key == 11'b10000110100) ? 46'b0100111110011001000110001101101111111001000001 :
(key == 11'b10000110101) ? 46'b0100111101111101100110101101101111010100111110 :
(key == 11'b10000110110) ? 46'b0100111101100010001000101101101110110000111111 :
(key == 11'b10000110111) ? 46'b0100111101000110101011101101101110001101000001 :
(key == 11'b10000111000) ? 46'b0100111100101011010000001101101101101001000111 :
(key == 11'b10000111001) ? 46'b0100111100001111110101001101101101000101001101 :
(key == 11'b10000111010) ? 46'b0100111011110100011011101101101100100001010111 :
(key == 11'b10000111011) ? 46'b0100111011011001000011001101101011111101100010 :
(key == 11'b10000111100) ? 46'b0100111010111101101011101101101011011001101111 :
(key == 11'b10000111101) ? 46'b0100111010100010010101101101101010110110000000 :
(key == 11'b10000111110) ? 46'b0100111010000111000000001101101010010010010001 :
(key == 11'b10000111111) ? 46'b0100111001101011101100001101101001101110100101 :
(key == 11'b10001000000) ? 46'b0100111001010000011001101101101001001010111100 :
(key == 11'b10001000001) ? 46'b0100111000110101000111101101101000100111010100 :
(key == 11'b10001000010) ? 46'b0100111000011001110111001101101000000011101111 :
(key == 11'b10001000011) ? 46'b0100110111111110100111101101100111100000001100 :
(key == 11'b10001000100) ? 46'b0100110111100011011001001101100110111100101011 :
(key == 11'b10001000101) ? 46'b0100110111001000001011101101100110011001001100 :
(key == 11'b10001000110) ? 46'b0100110110101100111111101101100101110101110000 :
(key == 11'b10001000111) ? 46'b0100110110010001110100001101100101010010010101 :
(key == 11'b10001001000) ? 46'b0100110101110110101010001101100100101110111101 :
(key == 11'b10001001001) ? 46'b0100110101011011100001001101100100001011100110 :
(key == 11'b10001001010) ? 46'b0100110101000000011001101101100011101000010011 :
(key == 11'b10001001011) ? 46'b0100110100100101010010101101100011000101000001 :
(key == 11'b10001001100) ? 46'b0100110100001010001101001101100010100001110001 :
(key == 11'b10001001101) ? 46'b0100110011101111001000101101100001111110100100 :
(key == 11'b10001001110) ? 46'b0100110011010100000101001101100001011011011000 :
(key == 11'b10001001111) ? 46'b0100110010111001000011001101100000111000001111 :
(key == 11'b10001010000) ? 46'b0100110010011110000001101101100000010101001000 :
(key == 11'b10001010001) ? 46'b0100110010000011000001101101011111110010000011 :
(key == 11'b10001010010) ? 46'b0100110001101000000010101101011111001111000000 :
(key == 11'b10001010011) ? 46'b0100110001001101000100101101011110101011111111 :
(key == 11'b10001010100) ? 46'b0100110000110010001000001101011110001001000001 :
(key == 11'b10001010101) ? 46'b0100110000010111001100001101011101100110000100 :
(key == 11'b10001010110) ? 46'b0100101111111100010001101101011101000011001010 :
(key == 11'b10001010111) ? 46'b0100101111100001011000001101011100100000010010 :
(key == 11'b10001011000) ? 46'b0100101111000110011111101101011011111101011100 :
(key == 11'b10001011001) ? 46'b0100101110101011101000001101011011011010101000 :
(key == 11'b10001011010) ? 46'b0100101110010000110001101101011010110111110110 :
(key == 11'b10001011011) ? 46'b0100101101110101111100101101011010010101000110 :
(key == 11'b10001011100) ? 46'b0100101101011011001000101101011001110010011001 :
(key == 11'b10001011101) ? 46'b0100101101000000010101101101011001001111101101 :
(key == 11'b10001011110) ? 46'b0100101100100101100011101101011000101101000100 :
(key == 11'b10001011111) ? 46'b0100101100001010110010101101011000001010011100 :
(key == 11'b10001100000) ? 46'b0100101011110000000010101101010111100111110111 :
(key == 11'b10001100001) ? 46'b0100101011010101010100001101010111000101010100 :
(key == 11'b10001100010) ? 46'b0100101010111010100110101101010110100010110011 :
(key == 11'b10001100011) ? 46'b0100101010011111111010001101010110000000010100 :
(key == 11'b10001100100) ? 46'b0100101010000101001110101101010101011101110111 :
(key == 11'b10001100101) ? 46'b0100101001101010100100001101010100111011011101 :
(key == 11'b10001100110) ? 46'b0100101001001111111010101101010100011001000100 :
(key == 11'b10001100111) ? 46'b0100101000110101010010101101010011110110101101 :
(key == 11'b10001101000) ? 46'b0100101000011010101011101101010011010100011001 :
(key == 11'b10001101001) ? 46'b0100101000000000000101001101010010110010000110 :
(key == 11'b10001101010) ? 46'b0100100111100101100000001101010010001111110110 :
(key == 11'b10001101011) ? 46'b0100100111001010111100001101010001101101100111 :
(key == 11'b10001101100) ? 46'b0100100110110000011001101101010001001011011100 :
(key == 11'b10001101101) ? 46'b0100100110010101110111101101010000101001010001 :
(key == 11'b10001101110) ? 46'b0100100101111011010110101101010000000111001001 :
(key == 11'b10001101111) ? 46'b0100100101100000110111001101001111100101000011 :
(key == 11'b10001110000) ? 46'b0100100101000110011000101101001111000010111111 :
(key == 11'b10001110001) ? 46'b0100100100101011111011001101001110100000111101 :
(key == 11'b10001110010) ? 46'b0100100100010001011110101101001101111110111101 :
(key == 11'b10001110011) ? 46'b0100100011110111000011001101001101011100111111 :
(key == 11'b10001110100) ? 46'b0100100011011100101000101101001100111011000011 :
(key == 11'b10001110101) ? 46'b0100100011000010001111001101001100011001001001 :
(key == 11'b10001110110) ? 46'b0100100010100111110111001101001011110111010010 :
(key == 11'b10001110111) ? 46'b0100100010001101011111101101001011010101011100 :
(key == 11'b10001111000) ? 46'b0100100001110011001001101101001010110011101000 :
(key == 11'b10001111001) ? 46'b0100100001011000110100101101001010010001110111 :
(key == 11'b10001111010) ? 46'b0100100000111110100000101101001001110000000111 :
(key == 11'b10001111011) ? 46'b0100100000100100001101101101001001001110011010 :
(key == 11'b10001111100) ? 46'b0100100000001001111011101101001000101100101110 :
(key == 11'b10001111101) ? 46'b0100011111101111101010101101001000001011000100 :
(key == 11'b10001111110) ? 46'b0100011111010101011011001101000111101001011101 :
(key == 11'b10001111111) ? 46'b0100011110111011001100001101000111000111110111 :
(key == 11'b10010000000) ? 46'b0100011110100000111110101101000110100110010100 :
(key == 11'b10010000001) ? 46'b0100011110000110110001101101000110000100110010 :
(key == 11'b10010000010) ? 46'b0100011101101100100110001101000101100011010011 :
(key == 11'b10010000011) ? 46'b0100011101010010011011101101000101000001110110 :
(key == 11'b10010000100) ? 46'b0100011100111000010010001101000100100000011010 :
(key == 11'b10010000101) ? 46'b0100011100011110001001101101000011111111000001 :
(key == 11'b10010000110) ? 46'b0100011100000100000010001101000011011101101001 :
(key == 11'b10010000111) ? 46'b0100011011101001111011101101000010111100010100 :
(key == 11'b10010001000) ? 46'b0100011011001111110110101101000010011011000001 :
(key == 11'b10010001001) ? 46'b0100011010110101110010001101000001111001101111 :
(key == 11'b10010001010) ? 46'b0100011010011011101110101101000001011000011111 :
(key == 11'b10010001011) ? 46'b0100011010000001101100101101000000110111010010 :
(key == 11'b10010001100) ? 46'b0100011001100111101011001101000000010110000110 :
(key == 11'b10010001101) ? 46'b0100011001001101101011001100111111110100111101 :
(key == 11'b10010001110) ? 46'b0100011000110011101100001100111111010011110101 :
(key == 11'b10010001111) ? 46'b0100011000011001101110001100111110110010110000 :
(key == 11'b10010010000) ? 46'b0100010111111111110000101100111110010001101100 :
(key == 11'b10010010001) ? 46'b0100010111100101110100101100111101110000101010 :
(key == 11'b10010010010) ? 46'b0100010111001011111001101100111101001111101011 :
(key == 11'b10010010011) ? 46'b0100010110110001111111101100111100101110101101 :
(key == 11'b10010010100) ? 46'b0100010110011000000111001100111100001101110010 :
(key == 11'b10010010101) ? 46'b0100010101111110001111001100111011101100111000 :
(key == 11'b10010010110) ? 46'b0100010101100100011000001100111011001100000000 :
(key == 11'b10010010111) ? 46'b0100010101001010100010001100111010101011001010 :
(key == 11'b10010011000) ? 46'b0100010100110000101101101100111010001010010111 :
(key == 11'b10010011001) ? 46'b0100010100010110111001101100111001101001100100 :
(key == 11'b10010011010) ? 46'b0100010011111101000110101100111001001000110100 :
(key == 11'b10010011011) ? 46'b0100010011100011010101001100111000101000000110 :
(key == 11'b10010011100) ? 46'b0100010011001001100100001100111000000111011010 :
(key == 11'b10010011101) ? 46'b0100010010101111110100101100110111100110110000 :
(key == 11'b10010011110) ? 46'b0100010010010110000101101100110111000110001000 :
(key == 11'b10010011111) ? 46'b0100010001111100011000001100110110100101100010 :
(key == 11'b10010100000) ? 46'b0100010001100010101011101100110110000100111101 :
(key == 11'b10010100001) ? 46'b0100010001001000111111101100110101100100011011 :
(key == 11'b10010100010) ? 46'b0100010000101111010101001100110101000011111010 :
(key == 11'b10010100011) ? 46'b0100010000010101101011101100110100100011011100 :
(key == 11'b10010100100) ? 46'b0100001111111100000011001100110100000010111111 :
(key == 11'b10010100101) ? 46'b0100001111100010011011101100110011100010100101 :
(key == 11'b10010100110) ? 46'b0100001111001000110100101100110011000010001100 :
(key == 11'b10010100111) ? 46'b0100001110101111001111001100110010100001110101 :
(key == 11'b10010101000) ? 46'b0100001110010101101010101100110010000001100000 :
(key == 11'b10010101001) ? 46'b0100001101111100000111001100110001100001001101 :
(key == 11'b10010101010) ? 46'b0100001101100010100100101100110001000000111100 :
(key == 11'b10010101011) ? 46'b0100001101001001000011001100110000100000101101 :
(key == 11'b10010101100) ? 46'b0100001100101111100010101100110000000000100000 :
(key == 11'b10010101101) ? 46'b0100001100010110000011001100101111100000010100 :
(key == 11'b10010101110) ? 46'b0100001011111100100100101100101111000000001011 :
(key == 11'b10010101111) ? 46'b0100001011100011000111001100101110100000000011 :
(key == 11'b10010110000) ? 46'b0100001011001001101010101100101101111111111101 :
(key == 11'b10010110001) ? 46'b0100001010110000001111001100101101011111111010 :
(key == 11'b10010110010) ? 46'b0100001010010110110100101100101100111111111000 :
(key == 11'b10010110011) ? 46'b0100001001111101011011001100101100011111111000 :
(key == 11'b10010110100) ? 46'b0100001001100100000010101100101011111111111010 :
(key == 11'b10010110101) ? 46'b0100001001001010101011001100101011011111111101 :
(key == 11'b10010110110) ? 46'b0100001000110001010100101100101011000000000011 :
(key == 11'b10010110111) ? 46'b0100001000010111111111001100101010100000001011 :
(key == 11'b10010111000) ? 46'b0100000111111110101010101100101010000000010100 :
(key == 11'b10010111001) ? 46'b0100000111100101010111001100101001100000011111 :
(key == 11'b10010111010) ? 46'b0100000111001100000100101100101001000000101101 :
(key == 11'b10010111011) ? 46'b0100000110110010110011001100101000100000111100 :
(key == 11'b10010111100) ? 46'b0100000110011001100010101100101000000001001101 :
(key == 11'b10010111101) ? 46'b0100000110000000010011001100100111100001011111 :
(key == 11'b10010111110) ? 46'b0100000101100111000100101100100111000001110100 :
(key == 11'b10010111111) ? 46'b0100000101001101110110101100100110100010001010 :
(key == 11'b10011000000) ? 46'b0100000100110100101010001100100110000010100011 :
(key == 11'b10011000001) ? 46'b0100000100011011011110101100100101100010111101 :
(key == 11'b10011000010) ? 46'b0100000100000010010100001100100101000011011001 :
(key == 11'b10011000011) ? 46'b0100000011101001001010101100100100100011110111 :
(key == 11'b10011000100) ? 46'b0100000011010000000001101100100100000100010111 :
(key == 11'b10011000101) ? 46'b0100000010110110111010001100100011100100111000 :
(key == 11'b10011000110) ? 46'b0100000010011101110011101100100011000101011100 :
(key == 11'b10011000111) ? 46'b0100000010000100101101101100100010100110000001 :
(key == 11'b10011001000) ? 46'b0100000001101011101001001100100010000110101001 :
(key == 11'b10011001001) ? 46'b0100000001010010100101101100100001100111010010 :
(key == 11'b10011001010) ? 46'b0100000000111001100010101100100001000111111100 :
(key == 11'b10011001011) ? 46'b0100000000100000100001001100100000101000101001 :
(key == 11'b10011001100) ? 46'b0100000000000111100000001100100000001001011000 :
(key == 11'b10011001101) ? 46'b0011111111101110100000001100011111101010001000 :
(key == 11'b10011001110) ? 46'b0011111111010101100001101100011111001010111010 :
(key == 11'b10011001111) ? 46'b0011111110111100100011101100011110101011101110 :
(key == 11'b10011010000) ? 46'b0011111110100011100110101100011110001100100100 :
(key == 11'b10011010001) ? 46'b0011111110001010101011001100011101101101011100 :
(key == 11'b10011010010) ? 46'b0011111101110001110000001100011101001110010110 :
(key == 11'b10011010011) ? 46'b0011111101011000110110001100011100101111010001 :
(key == 11'b10011010100) ? 46'b0011111100111111111101001100011100010000001110 :
(key == 11'b10011010101) ? 46'b0011111100100111000101001100011011110001001101 :
(key == 11'b10011010110) ? 46'b0011111100001110001110001100011011010010001110 :
(key == 11'b10011010111) ? 46'b0011111011110101010111101100011010110011010000 :
(key == 11'b10011011000) ? 46'b0011111011011100100010101100011010010100010100 :
(key == 11'b10011011001) ? 46'b0011111011000011101110101100011001110101011011 :
(key == 11'b10011011010) ? 46'b0011111010101010111011101100011001010110100011 :
(key == 11'b10011011011) ? 46'b0011111010010010001001001100011000110111101100 :
(key == 11'b10011011100) ? 46'b0011111001111001011000001100011000011000111000 :
(key == 11'b10011011101) ? 46'b0011111001100000100111101100010111111010000101 :
(key == 11'b10011011110) ? 46'b0011111001000111111000001100010111011011010100 :
(key == 11'b10011011111) ? 46'b0011111000101111001010001100010110111100100110 :
(key == 11'b10011100000) ? 46'b0011111000010110011100101100010110011101111000 :
(key == 11'b10011100001) ? 46'b0011110111111101110000001100010101111111001101 :
(key == 11'b10011100010) ? 46'b0011110111100101000100101100010101100000100011 :
(key == 11'b10011100011) ? 46'b0011110111001100011010001100010101000001111011 :
(key == 11'b10011100100) ? 46'b0011110110110011110000101100010100100011010101 :
(key == 11'b10011100101) ? 46'b0011110110011011000111101100010100000100110000 :
(key == 11'b10011100110) ? 46'b0011110110000010100000001100010011100110001110 :
(key == 11'b10011100111) ? 46'b0011110101101001111001101100010011000111101110 :
(key == 11'b10011101000) ? 46'b0011110101010001010011101100010010101001001110 :
(key == 11'b10011101001) ? 46'b0011110100111000101110101100010010001010110001 :
(key == 11'b10011101010) ? 46'b0011110100100000001011001100010001101100010110 :
(key == 11'b10011101011) ? 46'b0011110100000111101000001100010001001101111100 :
(key == 11'b10011101100) ? 46'b0011110011101111000110001100010000101111100100 :
(key == 11'b10011101101) ? 46'b0011110011010110100101001100010000010001001110 :
(key == 11'b10011101110) ? 46'b0011110010111110000101001100001111110010111001 :
(key == 11'b10011101111) ? 46'b0011110010100101100110001100001111010100100111 :
(key == 11'b10011110000) ? 46'b0011110010001101000111101100001110110110010110 :
(key == 11'b10011110001) ? 46'b0011110001110100101010101100001110011000000111 :
(key == 11'b10011110010) ? 46'b0011110001011100001110001100001101111001111001 :
(key == 11'b10011110011) ? 46'b0011110001000011110011001100001101011011101110 :
(key == 11'b10011110100) ? 46'b0011110000101011011000101100001100111101100100 :
(key == 11'b10011110101) ? 46'b0011110000010010111111001100001100011111011100 :
(key == 11'b10011110110) ? 46'b0011101111111010100110101100001100000001010101 :
(key == 11'b10011110111) ? 46'b0011101111100010001111001100001011100011010001 :
(key == 11'b10011111000) ? 46'b0011101111001001111000001100001011000101001101 :
(key == 11'b10011111001) ? 46'b0011101110110001100010101100001010100111001100 :
(key == 11'b10011111010) ? 46'b0011101110011001001101101100001010001001001100 :
(key == 11'b10011111011) ? 46'b0011101110000000111010001100001001101011001111 :
(key == 11'b10011111100) ? 46'b0011101101101000100111001100001001001101010011 :
(key == 11'b10011111101) ? 46'b0011101101010000010101001100001000101111011001 :
(key == 11'b10011111110) ? 46'b0011101100111000000100001100001000010001100000 :
(key == 11'b10011111111) ? 46'b0011101100011111110100001100000111110011101001 :
(key == 11'b10100000000) ? 46'b0011101100000111100101001100000111010101110100 :
(key == 11'b10100000001) ? 46'b0011101011101111010110101100000110111000000001 :
(key == 11'b10100000010) ? 46'b0011101011010111001001101100000110011010001111 :
(key == 11'b10100000011) ? 46'b0011101010111110111101001100000101111100011111 :
(key == 11'b10100000100) ? 46'b0011101010100110110001101100000101011110110001 :
(key == 11'b10100000101) ? 46'b0011101010001110100111001100000101000001000100 :
(key == 11'b10100000110) ? 46'b0011101001110110011101101100000100100011011010 :
(key == 11'b10100000111) ? 46'b0011101001011110010101001100000100000101110001 :
(key == 11'b10100001000) ? 46'b0011101001000110001101001100000011101000001001 :
(key == 11'b10100001001) ? 46'b0011101000101110000110101100000011001010100100 :
(key == 11'b10100001010) ? 46'b0011101000010110000000101100000010101100111111 :
(key == 11'b10100001011) ? 46'b0011100111111101111011101100000010001111011101 :
(key == 11'b10100001100) ? 46'b0011100111100101110111101100000001110001111101 :
(key == 11'b10100001101) ? 46'b0011100111001101110100101100000001010100011110 :
(key == 11'b10100001110) ? 46'b0011100110110101110010001100000000110111000000 :
(key == 11'b10100001111) ? 46'b0011100110011101110001001100000000011001100101 :
(key == 11'b10100010000) ? 46'b0011100110000101110000101011111111111100001011 :
(key == 11'b10100010001) ? 46'b0011100101101101110001001011111111011110110011 :
(key == 11'b10100010010) ? 46'b0011100101010101110010101011111111000001011100 :
(key == 11'b10100010011) ? 46'b0011100100111101110101001011111110100100001000 :
(key == 11'b10100010100) ? 46'b0011100100100101111000101011111110000110110101 :
(key == 11'b10100010101) ? 46'b0011100100001101111100101011111101101001100011 :
(key == 11'b10100010110) ? 46'b0011100011110110000010001011111101001100010100 :
(key == 11'b10100010111) ? 46'b0011100011011110001000001011111100101111000101 :
(key == 11'b10100011000) ? 46'b0011100011000110001111001011111100010001111001 :
(key == 11'b10100011001) ? 46'b0011100010101110010111001011111011110100101111 :
(key == 11'b10100011010) ? 46'b0011100010010110011111101011111011010111100101 :
(key == 11'b10100011011) ? 46'b0011100001111110101001101011111010111010011110 :
(key == 11'b10100011100) ? 46'b0011100001100110110100001011111010011101011000 :
(key == 11'b10100011101) ? 46'b0011100001001110111111101011111010000000010100 :
(key == 11'b10100011110) ? 46'b0011100000110111001100001011111001100011010010 :
(key == 11'b10100011111) ? 46'b0011100000011111011001101011111001000110010001 :
(key == 11'b10100100000) ? 46'b0011100000000111100111101011111000101001010010 :
(key == 11'b10100100001) ? 46'b0011011111101111110110101011111000001100010100 :
(key == 11'b10100100010) ? 46'b0011011111011000000111001011110111101111011001 :
(key == 11'b10100100011) ? 46'b0011011111000000010111101011110111010010011110 :
(key == 11'b10100100100) ? 46'b0011011110101000101001101011110110110101100110 :
(key == 11'b10100100101) ? 46'b0011011110010000111100101011110110011000101111 :
(key == 11'b10100100110) ? 46'b0011011101111001010000001011110101111011111010 :
(key == 11'b10100100111) ? 46'b0011011101100001100100101011110101011111000110 :
(key == 11'b10100101000) ? 46'b0011011101001001111010001011110101000010010101 :
(key == 11'b10100101001) ? 46'b0011011100110010010000101011110100100101100100 :
(key == 11'b10100101010) ? 46'b0011011100011010101000001011110100001000110110 :
(key == 11'b10100101011) ? 46'b0011011100000011000000001011110011101100001001 :
(key == 11'b10100101100) ? 46'b0011011011101011011001001011110011001111011101 :
(key == 11'b10100101101) ? 46'b0011011011010011110011001011110010110010110100 :
(key == 11'b10100101110) ? 46'b0011011010111100001110001011110010010110001100 :
(key == 11'b10100101111) ? 46'b0011011010100100101001101011110001111001100101 :
(key == 11'b10100110000) ? 46'b0011011010001101000110001011110001011101000000 :
(key == 11'b10100110001) ? 46'b0011011001110101100100001011110001000000011101 :
(key == 11'b10100110010) ? 46'b0011011001011110000010001011110000100011111011 :
(key == 11'b10100110011) ? 46'b0011011001000110100001101011110000000111011100 :
(key == 11'b10100110100) ? 46'b0011011000101111000010001011101111101010111110 :
(key == 11'b10100110101) ? 46'b0011011000010111100011001011101111001110100001 :
(key == 11'b10100110110) ? 46'b0011011000000000000101001011101110110010000110 :
(key == 11'b10100110111) ? 46'b0011010111101000100111101011101110010101101100 :
(key == 11'b10100111000) ? 46'b0011010111010001001011101011101101111001010100 :
(key == 11'b10100111001) ? 46'b0011010110111001110000001011101101011100111110 :
(key == 11'b10100111010) ? 46'b0011010110100010010101101011101101000000101001 :
(key == 11'b10100111011) ? 46'b0011010110001010111100001011101100100100010110 :
(key == 11'b10100111100) ? 46'b0011010101110011100011101011101100001000000101 :
(key == 11'b10100111101) ? 46'b0011010101011100001011101011101011101011110101 :
(key == 11'b10100111110) ? 46'b0011010101000100110100101011101011001111100110 :
(key == 11'b10100111111) ? 46'b0011010100101101011110101011101010110011011010 :
(key == 11'b10101000000) ? 46'b0011010100010110001001101011101010010111001111 :
(key == 11'b10101000001) ? 46'b0011010011111110110101001011101001111011000101 :
(key == 11'b10101000010) ? 46'b0011010011100111100010001011101001011110111110 :
(key == 11'b10101000011) ? 46'b0011010011010000001111001011101001000010110111 :
(key == 11'b10101000100) ? 46'b0011010010111000111101101011101000100110110010 :
(key == 11'b10101000101) ? 46'b0011010010100001101101001011101000001010110000 :
(key == 11'b10101000110) ? 46'b0011010010001010011101001011100111101110101110 :
(key == 11'b10101000111) ? 46'b0011010001110011001110001011100111010010101110 :
(key == 11'b10101001000) ? 46'b0011010001011011111111101011100110110110101111 :
(key == 11'b10101001001) ? 46'b0011010001000100110010101011100110011010110011 :
(key == 11'b10101001010) ? 46'b0011010000101101100110001011100101111110110111 :
(key == 11'b10101001011) ? 46'b0011010000010110011010101011100101100010111110 :
(key == 11'b10101001100) ? 46'b0011001111111111010000001011100101000111000110 :
(key == 11'b10101001101) ? 46'b0011001111101000000110001011100100101011001111 :
(key == 11'b10101001110) ? 46'b0011001111010000111101001011100100001111011010 :
(key == 11'b10101001111) ? 46'b0011001110111001110101001011100011110011100111 :
(key == 11'b10101010000) ? 46'b0011001110100010101110001011100011010111110101 :
(key == 11'b10101010001) ? 46'b0011001110001011100111101011100010111100000101 :
(key == 11'b10101010010) ? 46'b0011001101110100100010001011100010100000010110 :
(key == 11'b10101010011) ? 46'b0011001101011101011101101011100010000100101001 :
(key == 11'b10101010100) ? 46'b0011001101000110011010001011100001101000111110 :
(key == 11'b10101010101) ? 46'b0011001100101111010111001011100001001101010100 :
(key == 11'b10101010110) ? 46'b0011001100011000010101001011100000110001101011 :
(key == 11'b10101010111) ? 46'b0011001100000001010100001011100000010110000100 :
(key == 11'b10101011000) ? 46'b0011001011101010010011101011011111111010011111 :
(key == 11'b10101011001) ? 46'b0011001011010011010100101011011111011110111011 :
(key == 11'b10101011010) ? 46'b0011001010111100010110001011011111000011011001 :
(key == 11'b10101011011) ? 46'b0011001010100101011000001011011110100111111000 :
(key == 11'b10101011100) ? 46'b0011001010001110011011101011011110001100011001 :
(key == 11'b10101011101) ? 46'b0011001001110111011111101011011101110000111100 :
(key == 11'b10101011110) ? 46'b0011001001100000100100001011011101010101011111 :
(key == 11'b10101011111) ? 46'b0011001001001001101010001011011100111010000101 :
(key == 11'b10101100000) ? 46'b0011001000110010110000101011011100011110101100 :
(key == 11'b10101100001) ? 46'b0011001000011011111000001011011100000011010100 :
(key == 11'b10101100010) ? 46'b0011001000000101000000101011011011100111111111 :
(key == 11'b10101100011) ? 46'b0011000111101110001001101011011011001100101010 :
(key == 11'b10101100100) ? 46'b0011000111010111010011101011011010110001010111 :
(key == 11'b10101100101) ? 46'b0011000111000000011110101011011010010110000110 :
(key == 11'b10101100110) ? 46'b0011000110101001101010001011011001111010110110 :
(key == 11'b10101100111) ? 46'b0011000110010010110111001011011001011111101000 :
(key == 11'b10101101000) ? 46'b0011000101111100000100001011011001000100011011 :
(key == 11'b10101101001) ? 46'b0011000101100101010010101011011000101001010000 :
(key == 11'b10101101010) ? 46'b0011000101001110100001101011011000001110000110 :
(key == 11'b10101101011) ? 46'b0011000100110111110001101011010111110010111110 :
(key == 11'b10101101100) ? 46'b0011000100100001000010101011010111010111110111 :
(key == 11'b10101101101) ? 46'b0011000100001010010100001011010110111100110010 :
(key == 11'b10101101110) ? 46'b0011000011110011100110101011010110100001101110 :
(key == 11'b10101101111) ? 46'b0011000011011100111010001011010110000110101100 :
(key == 11'b10101110000) ? 46'b0011000011000110001110001011010101101011101011 :
(key == 11'b10101110001) ? 46'b0011000010101111100011101011010101010000101101 :
(key == 11'b10101110010) ? 46'b0011000010011000111001001011010100110101101111 :
(key == 11'b10101110011) ? 46'b0011000010000010010000001011010100011010110011 :
(key == 11'b10101110100) ? 46'b0011000001101011100111101011010011111111111000 :
(key == 11'b10101110101) ? 46'b0011000001010101000000001011010011100100111111 :
(key == 11'b10101110110) ? 46'b0011000000111110011001001011010011001010000111 :
(key == 11'b10101110111) ? 46'b0011000000100111110011101011010010101111010010 :
(key == 11'b10101111000) ? 46'b0011000000010001001110001011010010010100011100 :
(key == 11'b10101111001) ? 46'b0010111111111010101010001011010001111001101010 :
(key == 11'b10101111010) ? 46'b0010111111100100000110101011010001011110111000 :
(key == 11'b10101111011) ? 46'b0010111111001101100100001011010001000100001000 :
(key == 11'b10101111100) ? 46'b0010111110110111000010101011010000101001011001 :
(key == 11'b10101111101) ? 46'b0010111110100000100001101011010000001110101100 :
(key == 11'b10101111110) ? 46'b0010111110001010000001101011001111110100000000 :
(key == 11'b10101111111) ? 46'b0010111101110011100010101011001111011001010110 :
(key == 11'b10110000000) ? 46'b0010111101011101000100001011001110111110101101 :
(key == 11'b10110000001) ? 46'b0010111101000110100110101011001110100100000110 :
(key == 11'b10110000010) ? 46'b0010111100110000001001101011001110001001100000 :
(key == 11'b10110000011) ? 46'b0010111100011001101101101011001101101110111100 :
(key == 11'b10110000100) ? 46'b0010111100000011010010101011001101010100011001 :
(key == 11'b10110000101) ? 46'b0010111011101100111000101011001100111001111000 :
(key == 11'b10110000110) ? 46'b0010111011010110011111001011001100011111011000 :
(key == 11'b10110000111) ? 46'b0010111011000000000110101011001100000100111001 :
(key == 11'b10110001000) ? 46'b0010111010101001101111001011001011101010011101 :
(key == 11'b10110001001) ? 46'b0010111010010011011000001011001011010000000001 :
(key == 11'b10110001010) ? 46'b0010111001111101000010001011001010110101100111 :
(key == 11'b10110001011) ? 46'b0010111001100110101100101011001010011011001110 :
(key == 11'b10110001100) ? 46'b0010111001010000011000001011001010000000110111 :
(key == 11'b10110001101) ? 46'b0010111000111010000100101011001001100110100010 :
(key == 11'b10110001110) ? 46'b0010111000100011110001101011001001001100001101 :
(key == 11'b10110001111) ? 46'b0010111000001101011111101011001000110001111010 :
(key == 11'b10110010000) ? 46'b0010110111110111001110101011001000010111101001 :
(key == 11'b10110010001) ? 46'b0010110111100000111110001011000111111101011001 :
(key == 11'b10110010010) ? 46'b0010110111001010101110101011000111100011001011 :
(key == 11'b10110010011) ? 46'b0010110110110100100000001011000111001000111110 :
(key == 11'b10110010100) ? 46'b0010110110011110010010001011000110101110110011 :
(key == 11'b10110010101) ? 46'b0010110110001000000101001011000110010100101001 :
(key == 11'b10110010110) ? 46'b0010110101110001111001001011000101111010100000 :
(key == 11'b10110010111) ? 46'b0010110101011011101101101011000101100000011001 :
(key == 11'b10110011000) ? 46'b0010110101000101100011001011000101000110010011 :
(key == 11'b10110011001) ? 46'b0010110100101111011001001011000100101100001111 :
(key == 11'b10110011010) ? 46'b0010110100011001010000001011000100010010001100 :
(key == 11'b10110011011) ? 46'b0010110100000011001000001011000011111000001011 :
(key == 11'b10110011100) ? 46'b0010110011101101000000101011000011011110001011 :
(key == 11'b10110011101) ? 46'b0010110011010110111010001011000011000100001100 :
(key == 11'b10110011110) ? 46'b0010110011000000110100101011000010101010001111 :
(key == 11'b10110011111) ? 46'b0010110010101010101111101011000010010000010100 :
(key == 11'b10110100000) ? 46'b0010110010010100101011101011000001110110011001 :
(key == 11'b10110100001) ? 46'b0010110001111110101000001011000001011100100000 :
(key == 11'b10110100010) ? 46'b0010110001101000100101101011000001000010101001 :
(key == 11'b10110100011) ? 46'b0010110001010010100100001011000000101000110011 :
(key == 11'b10110100100) ? 46'b0010110000111100100011001011000000001110111110 :
(key == 11'b10110100101) ? 46'b0010110000100110100011001010111111110101001011 :
(key == 11'b10110100110) ? 46'b0010110000010000100011101010111111011011011001 :
(key == 11'b10110100111) ? 46'b0010101111111010100101001010111111000001101001 :
(key == 11'b10110101000) ? 46'b0010101111100100100111101010111110100111111010 :
(key == 11'b10110101001) ? 46'b0010101111001110101010101010111110001110001101 :
(key == 11'b10110101010) ? 46'b0010101110111000101110101010111101110100100001 :
(key == 11'b10110101011) ? 46'b0010101110100010110011101010111101011010110110 :
(key == 11'b10110101100) ? 46'b0010101110001100111001001010111101000001001101 :
(key == 11'b10110101101) ? 46'b0010101101110110111111101010111100100111100101 :
(key == 11'b10110101110) ? 46'b0010101101100001000110101010111100001101111111 :
(key == 11'b10110101111) ? 46'b0010101101001011001110101010111011110100011010 :
(key == 11'b10110110000) ? 46'b0010101100110101010111001010111011011010110110 :
(key == 11'b10110110001) ? 46'b0010101100011111100000101010111011000001010011 :
(key == 11'b10110110010) ? 46'b0010101100001001101011001010111010100111110011 :
(key == 11'b10110110011) ? 46'b0010101011110011110110101010111010001110010100 :
(key == 11'b10110110100) ? 46'b0010101011011110000010001010111001110100110101 :
(key == 11'b10110110101) ? 46'b0010101011001000001111001010111001011011011001 :
(key == 11'b10110110110) ? 46'b0010101010110010011100101010111001000001111101 :
(key == 11'b10110110111) ? 46'b0010101010011100101011001010111000101000100100 :
(key == 11'b10110111000) ? 46'b0010101010000110111010001010111000001111001011 :
(key == 11'b10110111001) ? 46'b0010101001110001001010001010110111110101110100 :
(key == 11'b10110111010) ? 46'b0010101001011011011010101010110111011100011110 :
(key == 11'b10110111011) ? 46'b0010101001000101101100001010110111000011001010 :
(key == 11'b10110111100) ? 46'b0010101000101111111110101010110110101001110111 :
(key == 11'b10110111101) ? 46'b0010101000011010010001101010110110010000100101 :
(key == 11'b10110111110) ? 46'b0010101000000100100101101010110101110111010101 :
(key == 11'b10110111111) ? 46'b0010100111101110111010001010110101011110000110 :
(key == 11'b10111000000) ? 46'b0010100111011001001111101010110101000100111001 :
(key == 11'b10111000001) ? 46'b0010100111000011100101101010110100101011101101 :
(key == 11'b10111000010) ? 46'b0010100110101101111100101010110100010010100010 :
(key == 11'b10111000011) ? 46'b0010100110011000010100101010110011111001011001 :
(key == 11'b10111000100) ? 46'b0010100110000010101101001010110011100000010001 :
(key == 11'b10111000101) ? 46'b0010100101101101000110101010110011000111001010 :
(key == 11'b10111000110) ? 46'b0010100101010111100000101010110010101110000101 :
(key == 11'b10111000111) ? 46'b0010100101000001111011101010110010010101000001 :
(key == 11'b10111001000) ? 46'b0010100100101100010111101010110001111011111111 :
(key == 11'b10111001001) ? 46'b0010100100010110110100001010110001100010111110 :
(key == 11'b10111001010) ? 46'b0010100100000001010001001010110001001001111110 :
(key == 11'b10111001011) ? 46'b0010100011101011101111101010110000110001000000 :
(key == 11'b10111001100) ? 46'b0010100011010110001110001010110000011000000010 :
(key == 11'b10111001101) ? 46'b0010100011000000101110001010101111111111000111 :
(key == 11'b10111001110) ? 46'b0010100010101011001110001010101111100110001100 :
(key == 11'b10111001111) ? 46'b0010100010010101101111101010101111001101010011 :
(key == 11'b10111010000) ? 46'b0010100010000000010001101010101110110100011100 :
(key == 11'b10111010001) ? 46'b0010100001101010110100001010101110011011100101 :
(key == 11'b10111010010) ? 46'b0010100001010101010111101010101110000010110000 :
(key == 11'b10111010011) ? 46'b0010100000111111111100001010101101101001111101 :
(key == 11'b10111010100) ? 46'b0010100000101010100001001010101101010001001011 :
(key == 11'b10111010101) ? 46'b0010100000010101000111001010101100111000011010 :
(key == 11'b10111010110) ? 46'b0010011111111111101101101010101100011111101010 :
(key == 11'b10111010111) ? 46'b0010011111101010010101001010101100000110111100 :
(key == 11'b10111011000) ? 46'b0010011111010100111101001010101011101110001111 :
(key == 11'b10111011001) ? 46'b0010011110111111100110001010101011010101100100 :
(key == 11'b10111011010) ? 46'b0010011110101010001111101010101010111100111001 :
(key == 11'b10111011011) ? 46'b0010011110010100111010001010101010100100010000 :
(key == 11'b10111011100) ? 46'b0010011101111111100101101010101010001011101001 :
(key == 11'b10111011101) ? 46'b0010011101101010010001101010101001110011000011 :
(key == 11'b10111011110) ? 46'b0010011101010100111110101010101001011010011110 :
(key == 11'b10111011111) ? 46'b0010011100111111101100001010101001000001111011 :
(key == 11'b10111100000) ? 46'b0010011100101010011010001010101000101001011000 :
(key == 11'b10111100001) ? 46'b0010011100010101001001001010101000010000110111 :
(key == 11'b10111100010) ? 46'b0010011011111111111001001010100111111000011000 :
(key == 11'b10111100011) ? 46'b0010011011101010101001101010100111011111111001 :
(key == 11'b10111100100) ? 46'b0010011011010101011011001010100111000111011100 :
(key == 11'b10111100101) ? 46'b0010011011000000001101001010100110101111000001 :
(key == 11'b10111100110) ? 46'b0010011010101011000000001010100110010110100110 :
(key == 11'b10111100111) ? 46'b0010011010010101110100001010100101111110001110 :
(key == 11'b10111101000) ? 46'b0010011010000000101000101010100101100101110110 :
(key == 11'b10111101001) ? 46'b0010011001101011011101101010100101001101100000 :
(key == 11'b10111101010) ? 46'b0010011001010110010011101010100100110101001011 :
(key == 11'b10111101011) ? 46'b0010011001000001001010001010100100011100110111 :
(key == 11'b10111101100) ? 46'b0010011000101100000001101010100100000100100100 :
(key == 11'b10111101101) ? 46'b0010011000010110111010001010100011101100010011 :
(key == 11'b10111101110) ? 46'b0010011000000001110011001010100011010100000100 :
(key == 11'b10111101111) ? 46'b0010010111101100101100101010100010111011110101 :
(key == 11'b10111110000) ? 46'b0010010111010111100111001010100010100011101000 :
(key == 11'b10111110001) ? 46'b0010010111000010100010101010100010001011011100 :
(key == 11'b10111110010) ? 46'b0010010110101101011110101010100001110011010001 :
(key == 11'b10111110011) ? 46'b0010010110011000011011001010100001011011001000 :
(key == 11'b10111110100) ? 46'b0010010110000011011000101010100001000011000000 :
(key == 11'b10111110101) ? 46'b0010010101101110010111001010100000101010111001 :
(key == 11'b10111110110) ? 46'b0010010101011001010110001010100000010010110100 :
(key == 11'b10111110111) ? 46'b0010010101000100010110001010011111111010110000 :
(key == 11'b10111111000) ? 46'b0010010100101111010110101010011111100010101101 :
(key == 11'b10111111001) ? 46'b0010010100011010010111101010011111001010101011 :
(key == 11'b10111111010) ? 46'b0010010100000101011001101010011110110010101011 :
(key == 11'b10111111011) ? 46'b0010010011110000011100101010011110011010101100 :
(key == 11'b10111111100) ? 46'b0010010011011011100000001010011110000010101111 :
(key == 11'b10111111101) ? 46'b0010010011000110100100101010011101101010110011 :
(key == 11'b10111111110) ? 46'b0010010010110001101001101010011101010010110111 :
(key == 11'b10111111111) ? 46'b0010010010011100101111001010011100111010111101 :
(key == 11'b11000000000) ? 46'b0010010010000111110101101010011100100011000101 :
(key == 11'b11000000001) ? 46'b0010010001110010111101001010011100001011001110 :
(key == 11'b11000000010) ? 46'b0010010001011110000101001010011011110011011000 :
(key == 11'b11000000011) ? 46'b0010010001001001001101101010011011011011100011 :
(key == 11'b11000000100) ? 46'b0010010000110100010111001010011011000011101111 :
(key == 11'b11000000101) ? 46'b0010010000011111100001101010011010101011111101 :
(key == 11'b11000000110) ? 46'b0010010000001010101100101010011010010100001100 :
(key == 11'b11000000111) ? 46'b0010001111110101111000001010011001111100011101 :
(key == 11'b11000001000) ? 46'b0010001111100001000100101010011001100100101110 :
(key == 11'b11000001001) ? 46'b0010001111001100010010001010011001001101000001 :
(key == 11'b11000001010) ? 46'b0010001110110111100000001010011000110101010110 :
(key == 11'b11000001011) ? 46'b0010001110100010101110101010011000011101101011 :
(key == 11'b11000001100) ? 46'b0010001110001101111110001010011000000110000010 :
(key == 11'b11000001101) ? 46'b0010001101111001001110001010010111101110011001 :
(key == 11'b11000001110) ? 46'b0010001101100100011111001010010111010110110011 :
(key == 11'b11000001111) ? 46'b0010001101001111110001001010010110111111001110 :
(key == 11'b11000010000) ? 46'b0010001100111011000011001010010110100111101001 :
(key == 11'b11000010001) ? 46'b0010001100100110010110101010010110010000000110 :
(key == 11'b11000010010) ? 46'b0010001100010001101010001010010101111000100100 :
(key == 11'b11000010011) ? 46'b0010001011111100111111001010010101100001000100 :
(key == 11'b11000010100) ? 46'b0010001011101000010100001010010101001001100101 :
(key == 11'b11000010101) ? 46'b0010001011010011101010001010010100110010000111 :
(key == 11'b11000010110) ? 46'b0010001010111111000001001010010100011010101010 :
(key == 11'b11000010111) ? 46'b0010001010101010011000101010010100000011001111 :
(key == 11'b11000011000) ? 46'b0010001010010101110001001010010011101011110101 :
(key == 11'b11000011001) ? 46'b0010001010000001001010001010010011010100011100 :
(key == 11'b11000011010) ? 46'b0010001001101100100011101010010010111101000100 :
(key == 11'b11000011011) ? 46'b0010001001010111111110001010010010100101101101 :
(key == 11'b11000011100) ? 46'b0010001001000011011001001010010010001110011000 :
(key == 11'b11000011101) ? 46'b0010001000101110110101001010010001110111000100 :
(key == 11'b11000011110) ? 46'b0010001000011010010001101010010001011111110001 :
(key == 11'b11000011111) ? 46'b0010001000000101101111001010010001001000011111 :
(key == 11'b11000100000) ? 46'b0010000111110001001101001010010000110001001111 :
(key == 11'b11000100001) ? 46'b0010000111011100101100001010010000011010000000 :
(key == 11'b11000100010) ? 46'b0010000111001000001011101010010000000010110010 :
(key == 11'b11000100011) ? 46'b0010000110110011101100001010001111101011100110 :
(key == 11'b11000100100) ? 46'b0010000110011111001101001010001111010100011010 :
(key == 11'b11000100101) ? 46'b0010000110001010101110101010001110111101010000 :
(key == 11'b11000100110) ? 46'b0010000101110110010001001010001110100110000111 :
(key == 11'b11000100111) ? 46'b0010000101100001110100001010001110001110111111 :
(key == 11'b11000101000) ? 46'b0010000101001101011000001010001101110111111001 :
(key == 11'b11000101001) ? 46'b0010000100111000111100101010001101100000110100 :
(key == 11'b11000101010) ? 46'b0010000100100100100010001010001101001001110000 :
(key == 11'b11000101011) ? 46'b0010000100010000001000001010001100110010101101 :
(key == 11'b11000101100) ? 46'b0010000011111011101111001010001100011011101011 :
(key == 11'b11000101101) ? 46'b0010000011100111010110101010001100000100101011 :
(key == 11'b11000101110) ? 46'b0010000011010010111110101010001011101101101100 :
(key == 11'b11000101111) ? 46'b0010000010111110100111101010001011010110101110 :
(key == 11'b11000110000) ? 46'b0010000010101010010001001010001010111111110001 :
(key == 11'b11000110001) ? 46'b0010000010010101111011101010001010101000110110 :
(key == 11'b11000110010) ? 46'b0010000010000001100110101010001010010001111011 :
(key == 11'b11000110011) ? 46'b0010000001101101010010101010001001111011000010 :
(key == 11'b11000110100) ? 46'b0010000001011000111111001010001001100100001010 :
(key == 11'b11000110101) ? 46'b0010000001000100101100001010001001001101010011 :
(key == 11'b11000110110) ? 46'b0010000000110000011010001010001000110110011110 :
(key == 11'b11000110111) ? 46'b0010000000011100001000101010001000011111101010 :
(key == 11'b11000111000) ? 46'b0010000000000111111000001010001000001000110111 :
(key == 11'b11000111001) ? 46'b0001111111110011101000001010000111110010000101 :
(key == 11'b11000111010) ? 46'b0001111111011111011001001010000111011011010100 :
(key == 11'b11000111011) ? 46'b0001111111001011001010101010000111000100100101 :
(key == 11'b11000111100) ? 46'b0001111110110110111100101010000110101101110110 :
(key == 11'b11000111101) ? 46'b0001111110100010101111101010000110010111001001 :
(key == 11'b11000111110) ? 46'b0001111110001110100011001010000110000000011101 :
(key == 11'b11000111111) ? 46'b0001111101111010010111101010000101101001110011 :
(key == 11'b11001000000) ? 46'b0001111101100110001100101010000101010011001001 :
(key == 11'b11001000001) ? 46'b0001111101010010000010101010000100111100100001 :
(key == 11'b11001000010) ? 46'b0001111100111101111001001010000100100101111010 :
(key == 11'b11001000011) ? 46'b0001111100101001110000001010000100001111010100 :
(key == 11'b11001000100) ? 46'b0001111100010101101000001010000011111000101111 :
(key == 11'b11001000101) ? 46'b0001111100000001100000101010000011100010001100 :
(key == 11'b11001000110) ? 46'b0001111011101101011001101010000011001011101001 :
(key == 11'b11001000111) ? 46'b0001111011011001010011101010000010110101001000 :
(key == 11'b11001001000) ? 46'b0001111011000101001110101010000010011110101000 :
(key == 11'b11001001001) ? 46'b0001111010110001001010001010000010001000001010 :
(key == 11'b11001001010) ? 46'b0001111010011101000110001010000001110001101100 :
(key == 11'b11001001011) ? 46'b0001111010001001000010101010000001011011001111 :
(key == 11'b11001001100) ? 46'b0001111001110101000000001010000001000100110100 :
(key == 11'b11001001101) ? 46'b0001111001100000111110101010000000101110011010 :
(key == 11'b11001001110) ? 46'b0001111001001100111101101010000000011000000001 :
(key == 11'b11001001111) ? 46'b0001111000111000111101001010000000000001101001 :
(key == 11'b11001010000) ? 46'b0001111000100100111101001001111111101011010010 :
(key == 11'b11001010001) ? 46'b0001111000010000111110001001111111010100111101 :
(key == 11'b11001010010) ? 46'b0001110111111101000000001001111110111110101001 :
(key == 11'b11001010011) ? 46'b0001110111101001000010001001111110101000010110 :
(key == 11'b11001010100) ? 46'b0001110111010101000101101001111110010010000100 :
(key == 11'b11001010101) ? 46'b0001110111000001001001001001111101111011110011 :
(key == 11'b11001010110) ? 46'b0001110110101101001101101001111101100101100100 :
(key == 11'b11001010111) ? 46'b0001110110011001010011001001111101001111010110 :
(key == 11'b11001011000) ? 46'b0001110110000101011000101001111100111001001000 :
(key == 11'b11001011001) ? 46'b0001110101110001011111001001111100100010111100 :
(key == 11'b11001011010) ? 46'b0001110101011101100110101001111100001100110001 :
(key == 11'b11001011011) ? 46'b0001110101001001101110101001111011110110100111 :
(key == 11'b11001011100) ? 46'b0001110100110101110111001001111011100000011111 :
(key == 11'b11001011101) ? 46'b0001110100100010000000101001111011001010010111 :
(key == 11'b11001011110) ? 46'b0001110100001110001010101001111010110100010001 :
(key == 11'b11001011111) ? 46'b0001110011111010010101001001111010011110001100 :
(key == 11'b11001100000) ? 46'b0001110011100110100000101001111010001000001000 :
(key == 11'b11001100001) ? 46'b0001110011010010101100101001111001110010000101 :
(key == 11'b11001100010) ? 46'b0001110010111110111001101001111001011100000011 :
(key == 11'b11001100011) ? 46'b0001110010101011000111001001111001000110000011 :
(key == 11'b11001100100) ? 46'b0001110010010111010101001001111000110000000011 :
(key == 11'b11001100101) ? 46'b0001110010000011100100001001111000011010000101 :
(key == 11'b11001100110) ? 46'b0001110001101111110011101001111000000100001000 :
(key == 11'b11001100111) ? 46'b0001110001011100000011101001110111101110001100 :
(key == 11'b11001101000) ? 46'b0001110001001000010100101001110111011000010001 :
(key == 11'b11001101001) ? 46'b0001110000110100100110001001110111000010010111 :
(key == 11'b11001101010) ? 46'b0001110000100000111000101001110110101100011111 :
(key == 11'b11001101011) ? 46'b0001110000001101001011101001110110010110100111 :
(key == 11'b11001101100) ? 46'b0001101111111001011111001001110110000000110001 :
(key == 11'b11001101101) ? 46'b0001101111100101110011001001110101101010111100 :
(key == 11'b11001101110) ? 46'b0001101111010010001000001001110101010101001000 :
(key == 11'b11001101111) ? 46'b0001101110111110011110001001110100111111010101 :
(key == 11'b11001110000) ? 46'b0001101110101010110100101001110100101001100011 :
(key == 11'b11001110001) ? 46'b0001101110010111001011101001110100010011110011 :
(key == 11'b11001110010) ? 46'b0001101110000011100011001001110011111110000011 :
(key == 11'b11001110011) ? 46'b0001101101101111111011101001110011101000010101 :
(key == 11'b11001110100) ? 46'b0001101101011100010100101001110011010010100111 :
(key == 11'b11001110101) ? 46'b0001101101001000101110101001110010111100111100 :
(key == 11'b11001110110) ? 46'b0001101100110101001000101001110010100111010000 :
(key == 11'b11001110111) ? 46'b0001101100100001100100001001110010010001100111 :
(key == 11'b11001111000) ? 46'b0001101100001101111111101001110001111011111110 :
(key == 11'b11001111001) ? 46'b0001101011111010011100001001110001100110010110 :
(key == 11'b11001111010) ? 46'b0001101011100110111001001001110001010000101111 :
(key == 11'b11001111011) ? 46'b0001101011010011010111001001110000111011001010 :
(key == 11'b11001111100) ? 46'b0001101010111111110101101001110000100101100110 :
(key == 11'b11001111101) ? 46'b0001101010101100010100101001110000010000000011 :
(key == 11'b11001111110) ? 46'b0001101010011000110100101001101111111010100001 :
(key == 11'b11001111111) ? 46'b0001101010000101010101001001101111100101000000 :
(key == 11'b11010000000) ? 46'b0001101001110001110110001001101111001111100000 :
(key == 11'b11010000001) ? 46'b0001101001011110011000001001101110111010000001 :
(key == 11'b11010000010) ? 46'b0001101001001010111010101001101110100100100100 :
(key == 11'b11010000011) ? 46'b0001101000110111011110001001101110001111001000 :
(key == 11'b11010000100) ? 46'b0001101000100100000001101001101101111001101100 :
(key == 11'b11010000101) ? 46'b0001101000010000100110001001101101100100010010 :
(key == 11'b11010000110) ? 46'b0001100111111101001011101001101101001110111001 :
(key == 11'b11010000111) ? 46'b0001100111101001110001001001101100111001100000 :
(key == 11'b11010001000) ? 46'b0001100111010110011000001001101100100100001010 :
(key == 11'b11010001001) ? 46'b0001100111000010111111001001101100001110110100 :
(key == 11'b11010001010) ? 46'b0001100110101111100111001001101011111001011111 :
(key == 11'b11010001011) ? 46'b0001100110011100001111101001101011100100001100 :
(key == 11'b11010001100) ? 46'b0001100110001000111000101001101011001110111001 :
(key == 11'b11010001101) ? 46'b0001100101110101100010101001101010111001100111 :
(key == 11'b11010001110) ? 46'b0001100101100010001101001001101010100100010111 :
(key == 11'b11010001111) ? 46'b0001100101001110111000001001101010001111001000 :
(key == 11'b11010010000) ? 46'b0001100100111011100100001001101001111001111010 :
(key == 11'b11010010001) ? 46'b0001100100101000010000101001101001100100101101 :
(key == 11'b11010010010) ? 46'b0001100100010100111101101001101001001111100000 :
(key == 11'b11010010011) ? 46'b0001100100000001101011101001101000111010010110 :
(key == 11'b11010010100) ? 46'b0001100011101110011010001001101000100101001100 :
(key == 11'b11010010101) ? 46'b0001100011011011001001001001101000010000000011 :
(key == 11'b11010010110) ? 46'b0001100011000111111001001001100111111010111011 :
(key == 11'b11010010111) ? 46'b0001100010110100101001101001100111100101110101 :
(key == 11'b11010011000) ? 46'b0001100010100001011010101001100111010000101111 :
(key == 11'b11010011001) ? 46'b0001100010001110001100101001100110111011101011 :
(key == 11'b11010011010) ? 46'b0001100001111010111111001001100110100110101000 :
(key == 11'b11010011011) ? 46'b0001100001100111110010001001100110010001100110 :
(key == 11'b11010011100) ? 46'b0001100001010100100110001001100101111100100101 :
(key == 11'b11010011101) ? 46'b0001100001000001011010101001100101100111100101 :
(key == 11'b11010011110) ? 46'b0001100000101110001111101001100101010010100110 :
(key == 11'b11010011111) ? 46'b0001100000011011000101001001100100111101100111 :
(key == 11'b11010100000) ? 46'b0001100000000111111011101001100100101000101011 :
(key == 11'b11010100001) ? 46'b0001011111110100110010101001100100010011101111 :
(key == 11'b11010100010) ? 46'b0001011111100001101010101001100011111110110101 :
(key == 11'b11010100011) ? 46'b0001011111001110100010101001100011101001111011 :
(key == 11'b11010100100) ? 46'b0001011110111011011011101001100011010101000010 :
(key == 11'b11010100101) ? 46'b0001011110101000010101101001100011000000001011 :
(key == 11'b11010100110) ? 46'b0001011110010101001111101001100010101011010100 :
(key == 11'b11010100111) ? 46'b0001011110000010001010101001100010010110011111 :
(key == 11'b11010101000) ? 46'b0001011101101111000110101001100010000001101011 :
(key == 11'b11010101001) ? 46'b0001011101011100000010101001100001101100110111 :
(key == 11'b11010101010) ? 46'b0001011101001000111111101001100001011000000101 :
(key == 11'b11010101011) ? 46'b0001011100110101111101001001100001000011010100 :
(key == 11'b11010101100) ? 46'b0001011100100010111011101001100000101110100101 :
(key == 11'b11010101101) ? 46'b0001011100001111111010001001100000011001110101 :
(key == 11'b11010101110) ? 46'b0001011011111100111001101001100000000101000111 :
(key == 11'b11010101111) ? 46'b0001011011101001111010001001011111110000011011 :
(key == 11'b11010110000) ? 46'b0001011011010110111010101001011111011011101111 :
(key == 11'b11010110001) ? 46'b0001011011000011111100001001011111000111000100 :
(key == 11'b11010110010) ? 46'b0001011010110000111110001001011110110010011010 :
(key == 11'b11010110011) ? 46'b0001011010011110000001001001011110011101110010 :
(key == 11'b11010110100) ? 46'b0001011010001011000100101001011110001001001010 :
(key == 11'b11010110101) ? 46'b0001011001111000001000101001011101110100100100 :
(key == 11'b11010110110) ? 46'b0001011001100101001101001001011101011111111110 :
(key == 11'b11010110111) ? 46'b0001011001010010010010101001011101001011011010 :
(key == 11'b11010111000) ? 46'b0001011000111111011000101001011100110110110111 :
(key == 11'b11010111001) ? 46'b0001011000101100011111001001011100100010010100 :
(key == 11'b11010111010) ? 46'b0001011000011001100110001001011100001101110011 :
(key == 11'b11010111011) ? 46'b0001011000000110101110001001011011111001010011 :
(key == 11'b11010111100) ? 46'b0001010111110011110110101001011011100100110011 :
(key == 11'b11010111101) ? 46'b0001010111100001000000001001011011010000010110 :
(key == 11'b11010111110) ? 46'b0001010111001110001001101001011010111011111000 :
(key == 11'b11010111111) ? 46'b0001010110111011010100001001011010100111011100 :
(key == 11'b11011000000) ? 46'b0001010110101000011111001001011010010011000001 :
(key == 11'b11011000001) ? 46'b0001010110010101101011001001011001111110100111 :
(key == 11'b11011000010) ? 46'b0001010110000010110111001001011001101010001110 :
(key == 11'b11011000011) ? 46'b0001010101110000000100001001011001010101110110 :
(key == 11'b11011000100) ? 46'b0001010101011101010010001001011001000001100000 :
(key == 11'b11011000101) ? 46'b0001010101001010100000001001011000101101001001 :
(key == 11'b11011000110) ? 46'b0001010100110111101111001001011000011000110101 :
(key == 11'b11011000111) ? 46'b0001010100100100111110101001011000000100100001 :
(key == 11'b11011001000) ? 46'b0001010100010010001110101001010111110000001110 :
(key == 11'b11011001001) ? 46'b0001010011111111011111101001010111011011111100 :
(key == 11'b11011001010) ? 46'b0001010011101100110001001001010111000111101100 :
(key == 11'b11011001011) ? 46'b0001010011011010000011001001010110110011011100 :
(key == 11'b11011001100) ? 46'b0001010011000111010110001001010110011111001110 :
(key == 11'b11011001101) ? 46'b0001010010110100101001001001010110001011000000 :
(key == 11'b11011001110) ? 46'b0001010010100001111101001001010101110110110011 :
(key == 11'b11011001111) ? 46'b0001010010001111010001101001010101100010101000 :
(key == 11'b11011010000) ? 46'b0001010001111100100111001001010101001110011101 :
(key == 11'b11011010001) ? 46'b0001010001101001111101001001010100111010010100 :
(key == 11'b11011010010) ? 46'b0001010001010111010011101001010100100110001011 :
(key == 11'b11011010011) ? 46'b0001010001000100101010101001010100010010000100 :
(key == 11'b11011010100) ? 46'b0001010000110010000010001001010011111101111101 :
(key == 11'b11011010101) ? 46'b0001010000011111011010101001010011101001111000 :
(key == 11'b11011010110) ? 46'b0001010000001100110011101001010011010101110011 :
(key == 11'b11011010111) ? 46'b0001001111111010001101001001010011000001110000 :
(key == 11'b11011011000) ? 46'b0001001111100111100111101001010010101101101110 :
(key == 11'b11011011001) ? 46'b0001001111010101000010101001010010011001101100 :
(key == 11'b11011011010) ? 46'b0001001111000010011110001001010010000101101100 :
(key == 11'b11011011011) ? 46'b0001001110101111111010001001010001110001101100 :
(key == 11'b11011011100) ? 46'b0001001110011101010110101001010001011101101110 :
(key == 11'b11011011101) ? 46'b0001001110001010110100001001010001001001110000 :
(key == 11'b11011011110) ? 46'b0001001101111000010010001001010000110101110100 :
(key == 11'b11011011111) ? 46'b0001001101100101110000101001010000100001111001 :
(key == 11'b11011100000) ? 46'b0001001101010011010000001001010000001101111110 :
(key == 11'b11011100001) ? 46'b0001001101000000110000001001001111111010000101 :
(key == 11'b11011100010) ? 46'b0001001100101110010000101001001111100110001101 :
(key == 11'b11011100011) ? 46'b0001001100011011110001101001001111010010010101 :
(key == 11'b11011100100) ? 46'b0001001100001001010011001001001110111110011111 :
(key == 11'b11011100101) ? 46'b0001001011110110110101101001001110101010101010 :
(key == 11'b11011100110) ? 46'b0001001011100100011000101001001110010110110101 :
(key == 11'b11011100111) ? 46'b0001001011010001111100001001001110000011000010 :
(key == 11'b11011101000) ? 46'b0001001010111111100000101001001101101111010000 :
(key == 11'b11011101001) ? 46'b0001001010101101000101001001001101011011011110 :
(key == 11'b11011101010) ? 46'b0001001010011010101010101001001101000111101110 :
(key == 11'b11011101011) ? 46'b0001001010001000010000101001001100110011111110 :
(key == 11'b11011101100) ? 46'b0001001001110101110111101001001100100000010000 :
(key == 11'b11011101101) ? 46'b0001001001100011011110101001001100001100100011 :
(key == 11'b11011101110) ? 46'b0001001001010001000110101001001011111000110110 :
(key == 11'b11011101111) ? 46'b0001001000111110101111001001001011100101001011 :
(key == 11'b11011110000) ? 46'b0001001000101100011000101001001011010001100001 :
(key == 11'b11011110001) ? 46'b0001001000011010000010001001001010111101110111 :
(key == 11'b11011110010) ? 46'b0001001000000111101100101001001010101010001111 :
(key == 11'b11011110011) ? 46'b0001000111110101010111101001001010010110100111 :
(key == 11'b11011110100) ? 46'b0001000111100011000011001001001010000011000001 :
(key == 11'b11011110101) ? 46'b0001000111010000101111001001001001101111011011 :
(key == 11'b11011110110) ? 46'b0001000110111110011100001001001001011011110111 :
(key == 11'b11011110111) ? 46'b0001000110101100001001101001001001001000010011 :
(key == 11'b11011111000) ? 46'b0001000110011001110111101001001000110100110001 :
(key == 11'b11011111001) ? 46'b0001000110000111100110001001001000100001001111 :
(key == 11'b11011111010) ? 46'b0001000101110101010101101001001000001101101111 :
(key == 11'b11011111011) ? 46'b0001000101100011000101101001000111111010001111 :
(key == 11'b11011111100) ? 46'b0001000101010000110110001001000111100110110000 :
(key == 11'b11011111101) ? 46'b0001000100111110100111001001000111010011010011 :
(key == 11'b11011111110) ? 46'b0001000100101100011000101001000110111111110110 :
(key == 11'b11011111111) ? 46'b0001000100011010001011001001000110101100011010 :
(key == 11'b11100000000) ? 46'b0001000100000111111110001001000110011001000000 :
(key == 11'b11100000001) ? 46'b0001000011110101110001101001000110000101100110 :
(key == 11'b11100000010) ? 46'b0001000011100011100101101001000101110010001101 :
(key == 11'b11100000011) ? 46'b0001000011010001011010001001000101011110110101 :
(key == 11'b11100000100) ? 46'b0001000010111111001111101001000101001011011110 :
(key == 11'b11100000101) ? 46'b0001000010101101000101101001000100111000001000 :
(key == 11'b11100000110) ? 46'b0001000010011010111100001001000100100100110011 :
(key == 11'b11100000111) ? 46'b0001000010001000110011001001000100010001011111 :
(key == 11'b11100001000) ? 46'b0001000001110110101011001001000011111110001100 :
(key == 11'b11100001001) ? 46'b0001000001100100100011101001000011101010111010 :
(key == 11'b11100001010) ? 46'b0001000001010010011100001001000011010111101001 :
(key == 11'b11100001011) ? 46'b0001000001000000010110001001000011000100011001 :
(key == 11'b11100001100) ? 46'b0001000000101110010000001001000010110001001010 :
(key == 11'b11100001101) ? 46'b0001000000011100001010101001000010011101111011 :
(key == 11'b11100001110) ? 46'b0001000000001010000110001001000010001010101110 :
(key == 11'b11100001111) ? 46'b0000111111111000000010001001000001110111100010 :
(key == 11'b11100010000) ? 46'b0000111111100101111110101001000001100100010110 :
(key == 11'b11100010001) ? 46'b0000111111010011111100001001000001010001001100 :
(key == 11'b11100010010) ? 46'b0000111111000001111001101001000000111110000011 :
(key == 11'b11100010011) ? 46'b0000111110101111111000001001000000101010111010 :
(key == 11'b11100010100) ? 46'b0000111110011101110111001001000000010111110011 :
(key == 11'b11100010101) ? 46'b0000111110001011110110101001000000000100101100 :
(key == 11'b11100010110) ? 46'b0000111101111001110110101000111111110001100110 :
(key == 11'b11100010111) ? 46'b0000111101100111110111101000111111011110100010 :
(key == 11'b11100011000) ? 46'b0000111101010101111000101000111111001011011110 :
(key == 11'b11100011001) ? 46'b0000111101000011111010101000111110111000011011 :
(key == 11'b11100011010) ? 46'b0000111100110001111101001000111110100101011001 :
(key == 11'b11100011011) ? 46'b0000111100100000000000101000111110010010011001 :
(key == 11'b11100011100) ? 46'b0000111100001110000100001000111101111111011000 :
(key == 11'b11100011101) ? 46'b0000111011111100001000101000111101101100011010 :
(key == 11'b11100011110) ? 46'b0000111011101010001101001000111101011001011011 :
(key == 11'b11100011111) ? 46'b0000111011011000010010101000111101000110011110 :
(key == 11'b11100100000) ? 46'b0000111011000110011001001000111100110011100010 :
(key == 11'b11100100001) ? 46'b0000111010110100011111101000111100100000100111 :
(key == 11'b11100100010) ? 46'b0000111010100010100111001000111100001101101101 :
(key == 11'b11100100011) ? 46'b0000111010010000101110101000111011111010110011 :
(key == 11'b11100100100) ? 46'b0000111001111110110111001000111011100111111010 :
(key == 11'b11100100101) ? 46'b0000111001101101000000001000111011010101000011 :
(key == 11'b11100100110) ? 46'b0000111001011011001010001000111011000010001101 :
(key == 11'b11100100111) ? 46'b0000111001001001010100001000111010101111010111 :
(key == 11'b11100101000) ? 46'b0000111000110111011111001000111010011100100010 :
(key == 11'b11100101001) ? 46'b0000111000100101101010001000111010001001101110 :
(key == 11'b11100101010) ? 46'b0000111000010011110110001000111001110110111011 :
(key == 11'b11100101011) ? 46'b0000111000000010000011001000111001100100001010 :
(key == 11'b11100101100) ? 46'b0000110111110000010000001000111001010001011001 :
(key == 11'b11100101101) ? 46'b0000110111011110011101101000111000111110101000 :
(key == 11'b11100101110) ? 46'b0000110111001100101100001000111000101011111001 :
(key == 11'b11100101111) ? 46'b0000110110111010111011001000111000011001001011 :
(key == 11'b11100110000) ? 46'b0000110110101001001010101000111000000110011110 :
(key == 11'b11100110001) ? 46'b0000110110010111011010101000110111110011110001 :
(key == 11'b11100110010) ? 46'b0000110110000101101011001000110111100001000110 :
(key == 11'b11100110011) ? 46'b0000110101110011111100101000110111001110011100 :
(key == 11'b11100110100) ? 46'b0000110101100010001110101000110110111011110010 :
(key == 11'b11100110101) ? 46'b0000110101010000100000101000110110101001001001 :
(key == 11'b11100110110) ? 46'b0000110100111110110011101000110110010110100001 :
(key == 11'b11100110111) ? 46'b0000110100101101000111101000110110000011111011 :
(key == 11'b11100111000) ? 46'b0000110100011011011011101000110101110001010101 :
(key == 11'b11100111001) ? 46'b0000110100001001110000101000110101011110110000 :
(key == 11'b11100111010) ? 46'b0000110011111000000101101000110101001100001011 :
(key == 11'b11100111011) ? 46'b0000110011100110011011101000110100111001101000 :
(key == 11'b11100111100) ? 46'b0000110011010100110010001000110100100111000110 :
(key == 11'b11100111101) ? 46'b0000110011000011001001001000110100010100100101 :
(key == 11'b11100111110) ? 46'b0000110010110001100000101000110100000010000100 :
(key == 11'b11100111111) ? 46'b0000110010011111111001001000110011101111100101 :
(key == 11'b11101000000) ? 46'b0000110010001110010001101000110011011101000110 :
(key == 11'b11101000001) ? 46'b0000110001111100101011001000110011001010101000 :
(key == 11'b11101000010) ? 46'b0000110001101011000101001000110010111000001011 :
(key == 11'b11101000011) ? 46'b0000110001011001011111101000110010100101110000 :
(key == 11'b11101000100) ? 46'b0000110001000111111010101000110010010011010100 :
(key == 11'b11101000101) ? 46'b0000110000110110010110101000110010000000111011 :
(key == 11'b11101000110) ? 46'b0000110000100100110010101000110001101110100001 :
(key == 11'b11101000111) ? 46'b0000110000010011001111101000110001011100001001 :
(key == 11'b11101001000) ? 46'b0000110000000001101101001000110001001001110010 :
(key == 11'b11101001001) ? 46'b0000101111110000001011001000110000110111011011 :
(key == 11'b11101001010) ? 46'b0000101111011110101001101000110000100101000110 :
(key == 11'b11101001011) ? 46'b0000101111001101001000101000110000010010110001 :
(key == 11'b11101001100) ? 46'b0000101110111011101000001000110000000000011101 :
(key == 11'b11101001101) ? 46'b0000101110101010001000101000101111101110001010 :
(key == 11'b11101001110) ? 46'b0000101110011000101001101000101111011011111000 :
(key == 11'b11101001111) ? 46'b0000101110000111001011001000101111001001100111 :
(key == 11'b11101010000) ? 46'b0000101101110101101101001000101110110111010111 :
(key == 11'b11101010001) ? 46'b0000101101100100001111101000101110100101001000 :
(key == 11'b11101010010) ? 46'b0000101101010010110010101000101110010010111001 :
(key == 11'b11101010011) ? 46'b0000101101000001010110001000101110000000101011 :
(key == 11'b11101010100) ? 46'b0000101100101111111010101000101101101110011111 :
(key == 11'b11101010101) ? 46'b0000101100011110011111001000101101011100010011 :
(key == 11'b11101010110) ? 46'b0000101100001101000100101000101101001010001000 :
(key == 11'b11101010111) ? 46'b0000101011111011101010101000101100110111111110 :
(key == 11'b11101011000) ? 46'b0000101011101010010001001000101100100101110101 :
(key == 11'b11101011001) ? 46'b0000101011011000111000001000101100010011101101 :
(key == 11'b11101011010) ? 46'b0000101011000111100000001000101100000001100110 :
(key == 11'b11101011011) ? 46'b0000101010110110001000001000101011101111011111 :
(key == 11'b11101011100) ? 46'b0000101010100100110001001000101011011101011010 :
(key == 11'b11101011101) ? 46'b0000101010010011011010101000101011001011010101 :
(key == 11'b11101011110) ? 46'b0000101010000010000100001000101010111001010001 :
(key == 11'b11101011111) ? 46'b0000101001110000101110101000101010100111001110 :
(key == 11'b11101100000) ? 46'b0000101001011111011010001000101010010101001101 :
(key == 11'b11101100001) ? 46'b0000101001001110000101101000101010000011001011 :
(key == 11'b11101100010) ? 46'b0000101000111100110001101000101001110001001011 :
(key == 11'b11101100011) ? 46'b0000101000101011011110101000101001011111001100 :
(key == 11'b11101100100) ? 46'b0000101000011010001011101000101001001101001101 :
(key == 11'b11101100101) ? 46'b0000101000001000111001101000101000111011001111 :
(key == 11'b11101100110) ? 46'b0000100111110111101000001000101000101001010011 :
(key == 11'b11101100111) ? 46'b0000100111100110010111001000101000010111010111 :
(key == 11'b11101101000) ? 46'b0000100111010101000110101000101000000101011100 :
(key == 11'b11101101001) ? 46'b0000100111000011110110101000100111110011100010 :
(key == 11'b11101101010) ? 46'b0000100110110010100111001000100111100001101000 :
(key == 11'b11101101011) ? 46'b0000100110100001011000101000100111001111110000 :
(key == 11'b11101101100) ? 46'b0000100110010000001010001000100110111101111000 :
(key == 11'b11101101101) ? 46'b0000100101111110111100101000100110101100000010 :
(key == 11'b11101101110) ? 46'b0000100101101101101111101000100110011010001100 :
(key == 11'b11101101111) ? 46'b0000100101011100100011001000100110001000010111 :
(key == 11'b11101110000) ? 46'b0000100101001011010111001000100101110110100011 :
(key == 11'b11101110001) ? 46'b0000100100111010001011101000100101100100110000 :
(key == 11'b11101110010) ? 46'b0000100100101001000000101000100101010010111101 :
(key == 11'b11101110011) ? 46'b0000100100010111110110101000100101000001001100 :
(key == 11'b11101110100) ? 46'b0000100100000110101100101000100100101111011011 :
(key == 11'b11101110101) ? 46'b0000100011110101100011101000100100011101101100 :
(key == 11'b11101110110) ? 46'b0000100011100100011010101000100100001011111100 :
(key == 11'b11101110111) ? 46'b0000100011010011010010101000100011111010001111 :
(key == 11'b11101111000) ? 46'b0000100011000010001011001000100011101000100001 :
(key == 11'b11101111001) ? 46'b0000100010110001000100001000100011010110110101 :
(key == 11'b11101111010) ? 46'b0000100010011111111101101000100011000101001010 :
(key == 11'b11101111011) ? 46'b0000100010001110111000001000100010110011011111 :
(key == 11'b11101111100) ? 46'b0000100001111101110010101000100010100001110101 :
(key == 11'b11101111101) ? 46'b0000100001101100101101101000100010010000001100 :
(key == 11'b11101111110) ? 46'b0000100001011011101001101000100001111110100101 :
(key == 11'b11101111111) ? 46'b0000100001001010100110001000100001101100111110 :
(key == 11'b11110000000) ? 46'b0000100000111001100010101000100001011011010111 :
(key == 11'b11110000001) ? 46'b0000100000101000100000001000100001001001110001 :
(key == 11'b11110000010) ? 46'b0000100000010111011110001000100000111000001101 :
(key == 11'b11110000011) ? 46'b0000100000000110011100101000100000100110101001 :
(key == 11'b11110000100) ? 46'b0000011111110101011011101000100000010101000110 :
(key == 11'b11110000101) ? 46'b0000011111100100011011001000100000000011100100 :
(key == 11'b11110000110) ? 46'b0000011111010011011011101000011111110010000011 :
(key == 11'b11110000111) ? 46'b0000011111000010011100001000011111100000100010 :
(key == 11'b11110001000) ? 46'b0000011110110001011101101000011111001111000011 :
(key == 11'b11110001001) ? 46'b0000011110100000011111001000011110111101100100 :
(key == 11'b11110001010) ? 46'b0000011110001111100001101000011110101100000110 :
(key == 11'b11110001011) ? 46'b0000011101111110100100101000011110011010101001 :
(key == 11'b11110001100) ? 46'b0000011101101101101000001000011110001001001101 :
(key == 11'b11110001101) ? 46'b0000011101011100101100001000011101110111110010 :
(key == 11'b11110001110) ? 46'b0000011101001011110000101000011101100110011000 :
(key == 11'b11110001111) ? 46'b0000011100111010110101101000011101010100111110 :
(key == 11'b11110010000) ? 46'b0000011100101001111011001000011101000011100101 :
(key == 11'b11110010001) ? 46'b0000011100011001000001001000011100110010001101 :
(key == 11'b11110010010) ? 46'b0000011100001000001000001000011100100000110110 :
(key == 11'b11110010011) ? 46'b0000011011110111001111001000011100001111011111 :
(key == 11'b11110010100) ? 46'b0000011011100110010111001000011011111110001010 :
(key == 11'b11110010101) ? 46'b0000011011010101011111101000011011101100110110 :
(key == 11'b11110010110) ? 46'b0000011011000100101000001000011011011011100001 :
(key == 11'b11110010111) ? 46'b0000011010110011110001101000011011001010001111 :
(key == 11'b11110011000) ? 46'b0000011010100010111011101000011010111000111100 :
(key == 11'b11110011001) ? 46'b0000011010010010000110001000011010100111101011 :
(key == 11'b11110011010) ? 46'b0000011010000001010001001000011010010110011011 :
(key == 11'b11110011011) ? 46'b0000011001110000011100101000011010000101001011 :
(key == 11'b11110011100) ? 46'b0000011001011111101000101000011001110011111100 :
(key == 11'b11110011101) ? 46'b0000011001001110110101101000011001100010101110 :
(key == 11'b11110011110) ? 46'b0000011000111110000010101000011001010001100001 :
(key == 11'b11110011111) ? 46'b0000011000101101010000001000011001000000010100 :
(key == 11'b11110100000) ? 46'b0000011000011100011110101000011000101111001001 :
(key == 11'b11110100001) ? 46'b0000011000001011101101101000011000011101111111 :
(key == 11'b11110100010) ? 46'b0000010111111010111100101000011000001100110101 :
(key == 11'b11110100011) ? 46'b0000010111101010001100101000010111111011101100 :
(key == 11'b11110100100) ? 46'b0000010111011001011101001000010111101010100100 :
(key == 11'b11110100101) ? 46'b0000010111001000101110001000010111011001011100 :
(key == 11'b11110100110) ? 46'b0000010110110111111111101000010111001000010110 :
(key == 11'b11110100111) ? 46'b0000010110100111010001101000010110110111010000 :
(key == 11'b11110101000) ? 46'b0000010110010110100100001000010110100110001011 :
(key == 11'b11110101001) ? 46'b0000010110000101110111001000010110010101000111 :
(key == 11'b11110101010) ? 46'b0000010101110101001010101000010110000100000011 :
(key == 11'b11110101011) ? 46'b0000010101100100011110101000010101110011000001 :
(key == 11'b11110101100) ? 46'b0000010101010011110011101000010101100001111111 :
(key == 11'b11110101101) ? 46'b0000010101000011001000101000010101010000111110 :
(key == 11'b11110101110) ? 46'b0000010100110010011110101000010100111111111110 :
(key == 11'b11110101111) ? 46'b0000010100100001110100101000010100101110111111 :
(key == 11'b11110110000) ? 46'b0000010100010001001011101000010100011110000001 :
(key == 11'b11110110001) ? 46'b0000010100000000100010101000010100001101000011 :
(key == 11'b11110110010) ? 46'b0000010011101111111010101000010011111100000110 :
(key == 11'b11110110011) ? 46'b0000010011011111010011001000010011101011001010 :
(key == 11'b11110110100) ? 46'b0000010011001110101100001000010011011010001111 :
(key == 11'b11110110101) ? 46'b0000010010111110000101101000010011001001010101 :
(key == 11'b11110110110) ? 46'b0000010010101101011111001000010010111000011011 :
(key == 11'b11110110111) ? 46'b0000010010011100111001101000010010100111100010 :
(key == 11'b11110111000) ? 46'b0000010010001100010101001000010010010110101011 :
(key == 11'b11110111001) ? 46'b0000010001111011110000101000010010000101110011 :
(key == 11'b11110111010) ? 46'b0000010001101011001100101000010001110100111101 :
(key == 11'b11110111011) ? 46'b0000010001011010101001001000010001100100000111 :
(key == 11'b11110111100) ? 46'b0000010001001010000110001000010001010011010010 :
(key == 11'b11110111101) ? 46'b0000010000111001100100001000010001000010011111 :
(key == 11'b11110111110) ? 46'b0000010000101001000010001000010000110001101011 :
(key == 11'b11110111111) ? 46'b0000010000011000100000101000010000100000111001 :
(key == 11'b11111000000) ? 46'b0000010000001000000000001000010000010000001000 :
(key == 11'b11111000001) ? 46'b0000001111110111011111101000001111111111010111 :
(key == 11'b11111000010) ? 46'b0000001111100111000000001000001111101110100111 :
(key == 11'b11111000011) ? 46'b0000001111010110100001001000001111011101111000 :
(key == 11'b11111000100) ? 46'b0000001111000110000010001000001111001101001001 :
(key == 11'b11111000101) ? 46'b0000001110110101100100001000001110111100011100 :
(key == 11'b11111000110) ? 46'b0000001110100101000110101000001110101011101111 :
(key == 11'b11111000111) ? 46'b0000001110010100101001001000001110011011000011 :
(key == 11'b11111001000) ? 46'b0000001110000100001100101000001110001010011000 :
(key == 11'b11111001001) ? 46'b0000001101110011110000101000001101111001101101 :
(key == 11'b11111001010) ? 46'b0000001101100011010101001000001101101001000100 :
(key == 11'b11111001011) ? 46'b0000001101010010111010001000001101011000011011 :
(key == 11'b11111001100) ? 46'b0000001101000010011111101000001101000111110011 :
(key == 11'b11111001101) ? 46'b0000001100110010000101101000001100110111001100 :
(key == 11'b11111001110) ? 46'b0000001100100001101100001000001100100110100101 :
(key == 11'b11111001111) ? 46'b0000001100010001010011001000001100010110000000 :
(key == 11'b11111010000) ? 46'b0000001100000000111010101000001100000101011011 :
(key == 11'b11111010001) ? 46'b0000001011110000100011001000001011110100110111 :
(key == 11'b11111010010) ? 46'b0000001011100000001011101000001011100100010100 :
(key == 11'b11111010011) ? 46'b0000001011001111110100101000001011010011110001 :
(key == 11'b11111010100) ? 46'b0000001010111111011110001000001011000011001111 :
(key == 11'b11111010101) ? 46'b0000001010101111001000101000001010110010101111 :
(key == 11'b11111010110) ? 46'b0000001010011110110011001000001010100010001110 :
(key == 11'b11111010111) ? 46'b0000001010001110011110001000001010010001101111 :
(key == 11'b11111011000) ? 46'b0000001001111110001010001000001010000001010000 :
(key == 11'b11111011001) ? 46'b0000001001101101110110001000001001110000110010 :
(key == 11'b11111011010) ? 46'b0000001001011101100011001000001001100000010110 :
(key == 11'b11111011011) ? 46'b0000001001001101010000001000001001001111111001 :
(key == 11'b11111011100) ? 46'b0000001000111100111110001000001000111111011110 :
(key == 11'b11111011101) ? 46'b0000001000101100101100001000001000101111000011 :
(key == 11'b11111011110) ? 46'b0000001000011100011011001000001000011110101001 :
(key == 11'b11111011111) ? 46'b0000001000001100001010001000001000001110010000 :
(key == 11'b11111100000) ? 46'b0000000111111011111010001000000111111101111000 :
(key == 11'b11111100001) ? 46'b0000000111101011101010101000000111101101100000 :
(key == 11'b11111100010) ? 46'b0000000111011011011011001000000111011101001001 :
(key == 11'b11111100011) ? 46'b0000000111001011001100101000000111001100110011 :
(key == 11'b11111100100) ? 46'b0000000110111010111110101000000110111100011110 :
(key == 11'b11111100101) ? 46'b0000000110101010110000101000000110101100001001 :
(key == 11'b11111100110) ? 46'b0000000110011010100011101000000110011011110101 :
(key == 11'b11111100111) ? 46'b0000000110001010010111001000000110001011100011 :
(key == 11'b11111101000) ? 46'b0000000101111010001011001000000101111011010000 :
(key == 11'b11111101001) ? 46'b0000000101101001111111101000000101101010111111 :
(key == 11'b11111101010) ? 46'b0000000101011001110100001000000101011010101110 :
(key == 11'b11111101011) ? 46'b0000000101001001101001101000000101001010011110 :
(key == 11'b11111101100) ? 46'b0000000100111001011111101000000100111010001111 :
(key == 11'b11111101101) ? 46'b0000000100101001010110001000000100101010000001 :
(key == 11'b11111101110) ? 46'b0000000100011001001101001000000100011001110011 :
(key == 11'b11111101111) ? 46'b0000000100001001000100101000000100001001100110 :
(key == 11'b11111110000) ? 46'b0000000011111000111100101000000011111001011010 :
(key == 11'b11111110001) ? 46'b0000000011101000110100101000000011101001001111 :
(key == 11'b11111110010) ? 46'b0000000011011000101101101000000011011001000100 :
(key == 11'b11111110011) ? 46'b0000000011001000100111001000000011001000111010 :
(key == 11'b11111110100) ? 46'b0000000010111000100001001000000010111000110001 :
(key == 11'b11111110101) ? 46'b0000000010101000011011101000000010101000101001 :
(key == 11'b11111110110) ? 46'b0000000010011000010110101000000010011000100001 :
(key == 11'b11111110111) ? 46'b0000000010001000010010001000000010001000011011 :
(key == 11'b11111111000) ? 46'b0000000001111000001110001000000001111000010101 :
(key == 11'b11111111001) ? 46'b0000000001101000001010101000000001101000001111 :
(key == 11'b11111111010) ? 46'b0000000001011000000111101000000001011000001011 :
(key == 11'b11111111011) ? 46'b0000000001001000000101001000000001001000000111 :
(key == 11'b11111111100) ? 46'b0000000000111000000011001000000000111000000100 :
(key == 11'b11111111101) ? 46'b0000000000101000000001101000000000101000000010 :
(key == 11'b11111111110) ? 46'b0000000000011000000000101000000000011000000000 :
(key == 11'b11111111111) ? 46'b0000000000001000000000001000000000001000000000 : 46'd0;


endmodule

`default_nettype wire
