`default_nettype none

module finv
   ( input wire [31:0] x,
     output wire [31:0] y,
     output wire ovf);

   /* TODO: assumptions
    * - inputs and output are not unnormal numbers or NaN or +-inf 
    * - if e is 0, the number is interpreted as +0
    * - overflow and underflow are treated as the same for ovf wire
    * - when underflow, y will be 0
    */

   // split sequence to each subsequence
   wire xs;
   wire [7:0] xe;
   wire [22:0] xm;
   assign {xs, xe, xm} = x;

   // calc s
   wire s;
   assign s = xs;

   // calc e
   wire [7:0] e;
   assign e = (xm == 23'd0) ? 8'd254 - xe : 8'd253 - xe; 

   // calc m
   wire [22:0] m;
   wire [45:0] val;
   wire [9:0] key;
   wire [12:0] v;
   assign {key, v} = xm;
   // lookup table and get constant and grad
   lookup_table lt(key, val);
   wire [23:0] constant;
   wire [24:0] grad;
   // constant supplements 1 at the MSB
   // grad supplements 00 at the LSB
   assign {constant, grad} = {1'b1, val, 2'b0};
   wire [37:0] tmp_grad; // 37 comes from 13 + 25 - 1
   assign tmp_grad = v * grad;
   wire [23:0] tmp_tmp_grad;
   // grad part is 14 bit long (meaning small)
   assign tmp_tmp_grad = {10'd0, tmp_grad[37:24]};
   wire [23:0] tmp_m;
   assign tmp_m = constant - tmp_tmp_grad;
   assign m = (xm == 23'd0) ? 23'd0 : tmp_m[22:0];

   assign y = {s, e, m};
   assign ovf = 0;

endmodule

module lookup_table
   ( input wire [9:0] key,
     output wire [45:0] value);

   assign value =
(key == 10'b0000000000) ? 46'b1111111111111111111110011111111100000000010100 :
(key == 10'b0000000001) ? 46'b1111111110000000000110011111110100000001110100 :
(key == 10'b0000000010) ? 46'b1111111100000000011110011111101100000100110011 :
(key == 10'b0000000011) ? 46'b1111111010000001000101111111100100001001010001 :
(key == 10'b0000000100) ? 46'b1111111000000001111101111111011100001111001111 :
(key == 10'b0000000101) ? 46'b1111110110000011000101011111010100010110101001 :
(key == 10'b0000000110) ? 46'b1111110100000100011100111111001100011111100011 :
(key == 10'b0000000111) ? 46'b1111110010000110000011111111000100101001111001 :
(key == 10'b0000001000) ? 46'b1111110000000111111010011110111100110101101101 :
(key == 10'b0000001001) ? 46'b1111101110001010000000011110110101000010111111 :
(key == 10'b0000001010) ? 46'b1111101100001100010110111110101101010001101100 :
(key == 10'b0000001011) ? 46'b1111101010001110111011111110100101100001110101 :
(key == 10'b0000001100) ? 46'b1111101000010001110000111110011101110011011100 :
(key == 10'b0000001101) ? 46'b1111100110010100110101011110010110000110011101 :
(key == 10'b0000001110) ? 46'b1111100100011000001001011110001110011010111001 :
(key == 10'b0000001111) ? 46'b1111100010011011101100011110000110110000110000 :
(key == 10'b0000010000) ? 46'b1111100000011111011110111101111111001000000001 :
(key == 10'b0000010001) ? 46'b1111011110100011100000111101110111100000101011 :
(key == 10'b0000010010) ? 46'b1111011100100111110001011101101111111010110001 :
(key == 10'b0000010011) ? 46'b1111011010101100010001111101101000010110001111 :
(key == 10'b0000010100) ? 46'b1111011000110001000000111101100000110011000110 :
(key == 10'b0000010101) ? 46'b1111010110110101111111011101011001010001010111 :
(key == 10'b0000010110) ? 46'b1111010100111011001101011101010001110000111111 :
(key == 10'b0000010111) ? 46'b1111010011000000101001011101001010010010000000 :
(key == 10'b0000011000) ? 46'b1111010001000110010100111101000010110100010110 :
(key == 10'b0000011001) ? 46'b1111001111001100001111011100111011011000000110 :
(key == 10'b0000011010) ? 46'b1111001101010010011000111100110011111101001100 :
(key == 10'b0000011011) ? 46'b1111001011011000110000011100101100100011101001 :
(key == 10'b0000011100) ? 46'b1111001001011111010111011100100101001011011101 :
(key == 10'b0000011101) ? 46'b1111000111100110001101011100011101110100100111 :
(key == 10'b0000011110) ? 46'b1111000101101101010001011100010110011111000101 :
(key == 10'b0000011111) ? 46'b1111000011110100100100111100001111001010111010 :
(key == 10'b0000100000) ? 46'b1111000001111100000110011100000111111000000100 :
(key == 10'b0000100001) ? 46'b1111000000000011110110111100000000100110100010 :
(key == 10'b0000100010) ? 46'b1110111110001011110101011011111001010110010101 :
(key == 10'b0000100011) ? 46'b1110111100010100000010111011110010000111011011 :
(key == 10'b0000100100) ? 46'b1110111010011100011110011011101010111001110110 :
(key == 10'b0000100101) ? 46'b1110111000100101001000111011100011101101100100 :
(key == 10'b0000100110) ? 46'b1110110110101110000001011011011100100010100100 :
(key == 10'b0000100111) ? 46'b1110110100110111000111111011010101011000111000 :
(key == 10'b0000101000) ? 46'b1110110011000000011101011011001110010000011111 :
(key == 10'b0000101001) ? 46'b1110110001001010000000111011000111001001010111 :
(key == 10'b0000101010) ? 46'b1110101111010011110010111011000000000011100010 :
(key == 10'b0000101011) ? 46'b1110101101011101110010011010111000111110111111 :
(key == 10'b0000101100) ? 46'b1110101011101000000000011010110001111011101100 :
(key == 10'b0000101101) ? 46'b1110101001110010011100011010101010111001101001 :
(key == 10'b0000101110) ? 46'b1110100111111101000110111010100011111000111001 :
(key == 10'b0000101111) ? 46'b1110100110000111111110111010011100111001011000 :
(key == 10'b0000110000) ? 46'b1110100100010011000101011010010101111011001001 :
(key == 10'b0000110001) ? 46'b1110100010011110011001011010001110111110001000 :
(key == 10'b0000110010) ? 46'b1110100000101001111011011010001000000010010110 :
(key == 10'b0000110011) ? 46'b1110011110110101101011111010000001000111110011 :
(key == 10'b0000110100) ? 46'b1110011101000001101001011001111010001110100001 :
(key == 10'b0000110101) ? 46'b1110011011001101110100111001110011010110011101 :
(key == 10'b0000110110) ? 46'b1110011001011010001101111001101100011111100110 :
(key == 10'b0000110111) ? 46'b1110010111100110110101011001100101101001111110 :
(key == 10'b0000111000) ? 46'b1110010101110011101001111001011110110101100100 :
(key == 10'b0000111001) ? 46'b1110010100000000101100011001011000000010010110 :
(key == 10'b0000111010) ? 46'b1110010010001101111011111001010001010000010101 :
(key == 10'b0000111011) ? 46'b1110010000011011011001011001001010011111100011 :
(key == 10'b0000111100) ? 46'b1110001110101001000100111001000011101111111100 :
(key == 10'b0000111101) ? 46'b1110001100110110111100111000111101000001100011 :
(key == 10'b0000111110) ? 46'b1110001011000101000010111000110110010100010100 :
(key == 10'b0000111111) ? 46'b1110001001010011010110011000101111101000010001 :
(key == 10'b0001000000) ? 46'b1110000111100001110111011000101000111101011011 :
(key == 10'b0001000001) ? 46'b1110000101110000100100111000100010010011101110 :
(key == 10'b0001000010) ? 46'b1110000011111111100000011000011011101011001111 :
(key == 10'b0001000011) ? 46'b1110000010001110101001011000010101000011111000 :
(key == 10'b0001000100) ? 46'b1110000000011101111111011000001110011101101100 :
(key == 10'b0001000101) ? 46'b1101111110101101100010011000000111111000101010 :
(key == 10'b0001000110) ? 46'b1101111100111101010010111000000001010100110011 :
(key == 10'b0001000111) ? 46'b1101111011001101001111110111111010110010000101 :
(key == 10'b0001001000) ? 46'b1101111001011101011001110111110100010000100000 :
(key == 10'b0001001001) ? 46'b1101110111101101110001010111101101110000000100 :
(key == 10'b0001001010) ? 46'b1101110101111110010101110111100111010000110001 :
(key == 10'b0001001011) ? 46'b1101110100001111000111110111100000110010100100 :
(key == 10'b0001001100) ? 46'b1101110010100000000101110111011010010101100010 :
(key == 10'b0001001101) ? 46'b1101110000110001010001010111010011111001101000 :
(key == 10'b0001001110) ? 46'b1101101111000010101001110111001101011110110101 :
(key == 10'b0001001111) ? 46'b1101101101010100001110110111000111000101001010 :
(key == 10'b0001010000) ? 46'b1101101011100110000000110111000000101100100101 :
(key == 10'b0001010001) ? 46'b1101101001110111111111010110111010010101000111 :
(key == 10'b0001010010) ? 46'b1101101000001010001010010110110011111110110010 :
(key == 10'b0001010011) ? 46'b1101100110011100100010010110101101101001100000 :
(key == 10'b0001010100) ? 46'b1101100100101111000111010110100111010101010110 :
(key == 10'b0001010101) ? 46'b1101100011000001111000110110100001000010010011 :
(key == 10'b0001010110) ? 46'b1101100001010100110110110110011010110000010100 :
(key == 10'b0001010111) ? 46'b1101011111101000000000110110010100011111011100 :
(key == 10'b0001011000) ? 46'b1101011101111011010111110110001110001111100111 :
(key == 10'b0001011001) ? 46'b1101011100001110111011110110001000000000111001 :
(key == 10'b0001011010) ? 46'b1101011010100010101011010110000001110011001101 :
(key == 10'b0001011011) ? 46'b1101011000110110100111110101111011100110100111 :
(key == 10'b0001011100) ? 46'b1101010111001010110000110101110101011011000101 :
(key == 10'b0001011101) ? 46'b1101010101011111000101110101101111010000101000 :
(key == 10'b0001011110) ? 46'b1101010011110011100111110101101001000111001101 :
(key == 10'b0001011111) ? 46'b1101010010001000010101010101100010111110110111 :
(key == 10'b0001100000) ? 46'b1101010000011101001111010101011100110111100011 :
(key == 10'b0001100001) ? 46'b1101001110110010010101010101010110110001010011 :
(key == 10'b0001100010) ? 46'b1101001101000111101000010101010000101100000101 :
(key == 10'b0001100011) ? 46'b1101001011011101000110110101001010100111111001 :
(key == 10'b0001100100) ? 46'b1101001001110010110001110101000100100100110000 :
(key == 10'b0001100101) ? 46'b1101001000001000101000010100111110100010101001 :
(key == 10'b0001100110) ? 46'b1101000110011110101011010100111000100001100100 :
(key == 10'b0001100111) ? 46'b1101000100110100111001110100110010100001100001 :
(key == 10'b0001101000) ? 46'b1101000011001011010101010100101100100010011101 :
(key == 10'b0001101001) ? 46'b1101000001100001111100010100100110100100011100 :
(key == 10'b0001101010) ? 46'b1100111111111000101110110100100000100111011100 :
(key == 10'b0001101011) ? 46'b1100111110001111101101110100011010101011011011 :
(key == 10'b0001101100) ? 46'b1100111100100110111000010100010100110000011011 :
(key == 10'b0001101101) ? 46'b1100111010111110001110110100001110110110011100 :
(key == 10'b0001101110) ? 46'b1100111001010101110000110100001000111101011110 :
(key == 10'b0001101111) ? 46'b1100110111101101011111010100000011000101011101 :
(key == 10'b0001110000) ? 46'b1100110110000101011001010011111101001110011101 :
(key == 10'b0001110001) ? 46'b1100110100011101011110110011110111011000011101 :
(key == 10'b0001110010) ? 46'b1100110010110101101111110011110001100011011011 :
(key == 10'b0001110011) ? 46'b1100110001001110001100110011101011101111010111 :
(key == 10'b0001110100) ? 46'b1100101111100110110101010011100101111100010011 :
(key == 10'b0001110101) ? 46'b1100101101111111101001010011100000001010001101 :
(key == 10'b0001110110) ? 46'b1100101100011000101001010011011010011001000110 :
(key == 10'b0001110111) ? 46'b1100101010110001110100010011010100101000111010 :
(key == 10'b0001111000) ? 46'b1100101001001011001011010011001110111001101110 :
(key == 10'b0001111001) ? 46'b1100100111100100101101010011001001001011011111 :
(key == 10'b0001111010) ? 46'b1100100101111110011010110011000011011110001111 :
(key == 10'b0001111011) ? 46'b1100100100011000010011110010111101110001111001 :
(key == 10'b0001111100) ? 46'b1100100010110010011000010010111000000110100011 :
(key == 10'b0001111101) ? 46'b1100100001001100101000010010110010011100001001 :
(key == 10'b0001111110) ? 46'b1100011111100111000011010010101100110010101001 :
(key == 10'b0001111111) ? 46'b1100011110000001101001110010100111001010000111 :
(key == 10'b0010000000) ? 46'b1100011100011100011011010010100001100010100010 :
(key == 10'b0010000001) ? 46'b1100011010110111011000010010011011111011110111 :
(key == 10'b0010000010) ? 46'b1100011001010010100000010010010110010110001000 :
(key == 10'b0010000011) ? 46'b1100010111101101110011110010010000110001010101 :
(key == 10'b0010000100) ? 46'b1100010110001001010001110010001011001101011101 :
(key == 10'b0010000101) ? 46'b1100010100100100111011110010000101101010100000 :
(key == 10'b0010000110) ? 46'b1100010011000000110000110010000000001000011111 :
(key == 10'b0010000111) ? 46'b1100010001011100110000010001111010100111010110 :
(key == 10'b0010001000) ? 46'b1100001111111000111010110001110101000111001010 :
(key == 10'b0010001001) ? 46'b1100001110010101010000110001101111100111110110 :
(key == 10'b0010001010) ? 46'b1100001100110001110001110001101010001001011110 :
(key == 10'b0010001011) ? 46'b1100001011001110011101010001100100101011111110 :
(key == 10'b0010001100) ? 46'b1100001001101011010011110001011111001111011000 :
(key == 10'b0010001101) ? 46'b1100001000001000010101010001011001110011101100 :
(key == 10'b0010001110) ? 46'b1100000110100101100001110001010100011000111010 :
(key == 10'b0010001111) ? 46'b1100000101000010111000110001001110111111000000 :
(key == 10'b0010010000) ? 46'b1100000011100000011011010001001001100101111111 :
(key == 10'b0010010001) ? 46'b1100000001111110000111110001000100001101110110 :
(key == 10'b0010010010) ? 46'b1100000000011011111111010000111110110110100110 :
(key == 10'b0010010011) ? 46'b1011111110111010000001110000111001100000001101 :
(key == 10'b0010010100) ? 46'b1011111101011000001110110000110100001010101110 :
(key == 10'b0010010101) ? 46'b1011111011110110100110010000101110110110000110 :
(key == 10'b0010010110) ? 46'b1011111010010101001000110000101001100010010101 :
(key == 10'b0010010111) ? 46'b1011111000110011110101110000100100001111011101 :
(key == 10'b0010011000) ? 46'b1011110111010010101101010000011110111101011011 :
(key == 10'b0010011001) ? 46'b1011110101110001101111010000011001101100010001 :
(key == 10'b0010011010) ? 46'b1011110100010000111011110000010100011011111110 :
(key == 10'b0010011011) ? 46'b1011110010110000010010110000001111001100100001 :
(key == 10'b0010011100) ? 46'b1011110001001111110100010000001001111101111010 :
(key == 10'b0010011101) ? 46'b1011101111101111100000110000000100110000001011 :
(key == 10'b0010011110) ? 46'b1011101110001111010111001111111111100011010000 :
(key == 10'b0010011111) ? 46'b1011101100101111010111101111111010010111001100 :
(key == 10'b0010100000) ? 46'b1011101011001111100011001111110101001011111110 :
(key == 10'b0010100001) ? 46'b1011101001101111111000101111110000000001100111 :
(key == 10'b0010100010) ? 46'b1011101000010000011000101111101010111000000011 :
(key == 10'b0010100011) ? 46'b1011100110110001000011001111100101101111010110 :
(key == 10'b0010100100) ? 46'b1011100101010001110111101111100000100111011101 :
(key == 10'b0010100101) ? 46'b1011100011110010110110001111011011100000011010 :
(key == 10'b0010100110) ? 46'b1011100010010011111111001111010110011010001010 :
(key == 10'b0010100111) ? 46'b1011100000110101010010101111010001010100110001 :
(key == 10'b0010101000) ? 46'b1011011111010110101111101111001100010000001001 :
(key == 10'b0010101001) ? 46'b1011011101111000010111001111000111001100011001 :
(key == 10'b0010101010) ? 46'b1011011100011010001001001111000010001001011010 :
(key == 10'b0010101011) ? 46'b1011011010111100000100101110111101000111010000 :
(key == 10'b0010101100) ? 46'b1011011001011110001010101110111000000101111010 :
(key == 10'b0010101101) ? 46'b1011011000000000011010101110110011000101011000 :
(key == 10'b0010101110) ? 46'b1011010110100010110100001110101110000101100111 :
(key == 10'b0010101111) ? 46'b1011010101000101010111101110101001000110101011 :
(key == 10'b0010110000) ? 46'b1011010011101000000101101110100100001000100001 :
(key == 10'b0010110001) ? 46'b1011010010001010111101101110011111001011001100 :
(key == 10'b0010110010) ? 46'b1011010000101101111111001110011010001110100111 :
(key == 10'b0010110011) ? 46'b1011001111010001001010101110010101010010110110 :
(key == 10'b0010110100) ? 46'b1011001101110100100000001110010000010111111000 :
(key == 10'b0010110101) ? 46'b1011001100010111111111101110001011011101101010 :
(key == 10'b0010110110) ? 46'b1011001010111011101000101110000110100100001111 :
(key == 10'b0010110111) ? 46'b1011001001011111011011101110000001101011100101 :
(key == 10'b0010111000) ? 46'b1011001000000011011000001101111100110011101110 :
(key == 10'b0010111001) ? 46'b1011000110100111011110101101110111111100101001 :
(key == 10'b0010111010) ? 46'b1011000101001011101110101101110011000110010100 :
(key == 10'b0010111011) ? 46'b1011000011110000001000001101101110010000110000 :
(key == 10'b0010111100) ? 46'b1011000010010100101011101101101001011011111110 :
(key == 10'b0010111101) ? 46'b1011000000111001011000101101100100100111111101 :
(key == 10'b0010111110) ? 46'b1010111111011110001111101101011111110100101100 :
(key == 10'b0010111111) ? 46'b1010111110000011001111101101011011000010001011 :
(key == 10'b0011000000) ? 46'b1010111100101000011001101101010110010000011010 :
(key == 10'b0011000001) ? 46'b1010111011001101101101001101010001011111011011 :
(key == 10'b0011000010) ? 46'b1010111001110011001010001101001100101111001010 :
(key == 10'b0011000011) ? 46'b1010111000011000110001001101000111111111101010 :
(key == 10'b0011000100) ? 46'b1010110110111110100001001101000011010000111001 :
(key == 10'b0011000101) ? 46'b1010110101100100011010001100111110100010111010 :
(key == 10'b0011000110) ? 46'b1010110100001010011101001100111001110101101000 :
(key == 10'b0011000111) ? 46'b1010110010110000101001101100110101001001000110 :
(key == 10'b0011001000) ? 46'b1010110001010110111111101100110000011101010011 :
(key == 10'b0011001001) ? 46'b1010101111111101011110101100101011110010001110 :
(key == 10'b0011001010) ? 46'b1010101110100100000110101100100111000111111011 :
(key == 10'b0011001011) ? 46'b1010101101001010111000101100100010011110010011 :
(key == 10'b0011001100) ? 46'b1010101011110001110011101100011101110101011100 :
(key == 10'b0011001101) ? 46'b1010101010011000111000001100011001001101010010 :
(key == 10'b0011001110) ? 46'b1010101001000000000101101100010100100101110110 :
(key == 10'b0011001111) ? 46'b1010100111100111011100101100001111111111001001 :
(key == 10'b0011010000) ? 46'b1010100110001110111100101100001011011001001001 :
(key == 10'b0011010001) ? 46'b1010100100110110100101101100000110110011110111 :
(key == 10'b0011010010) ? 46'b1010100011011110011000001100000010001111010011 :
(key == 10'b0011010011) ? 46'b1010100010000110010011101011111101101011011100 :
(key == 10'b0011010100) ? 46'b1010100000101110011000001011111001001000010010 :
(key == 10'b0011010101) ? 46'b1010011111010110100110001011110100100101110110 :
(key == 10'b0011010110) ? 46'b1010011101111110111100101011110000000100001000 :
(key == 10'b0011010111) ? 46'b1010011100100111011100101011101011100011000100 :
(key == 10'b0011011000) ? 46'b1010011011010000000101101011100111000010101110 :
(key == 10'b0011011001) ? 46'b1010011001111000110111101011100010100011000101 :
(key == 10'b0011011010) ? 46'b1010011000100001110010001011011110000100001001 :
(key == 10'b0011011011) ? 46'b1010010111001010110110101011011001100101110111 :
(key == 10'b0011011100) ? 46'b1010010101110100000011001011010101001000010100 :
(key == 10'b0011011101) ? 46'b1010010100011101011001001011010000101011011011 :
(key == 10'b0011011110) ? 46'b1010010011000110110111001011001100001111010000 :
(key == 10'b0011011111) ? 46'b1010010001110000011111001011000111110011101101 :
(key == 10'b0011100000) ? 46'b1010010000011010001111001011000011011000111001 :
(key == 10'b0011100001) ? 46'b1010001111000100001000101010111110111110101111 :
(key == 10'b0011100010) ? 46'b1010001101101110001010101010111010100101010001 :
(key == 10'b0011100011) ? 46'b1010001100011000010101101010110110001100011110 :
(key == 10'b0011100100) ? 46'b1010001011000010101001001010110001110100010110 :
(key == 10'b0011100101) ? 46'b1010001001101101000101101010101101011100111000 :
(key == 10'b0011100110) ? 46'b1010001000010111101010101010101001000110000110 :
(key == 10'b0011100111) ? 46'b1010000111000010011000001010100100101111111101 :
(key == 10'b0011101000) ? 46'b1010000101101101001110101010100000011010100000 :
(key == 10'b0011101001) ? 46'b1010000100011000001110001010011100000101101101 :
(key == 10'b0011101010) ? 46'b1010000011000011010101101010010111110001100100 :
(key == 10'b0011101011) ? 46'b1010000001101110100110001010010011011110000110 :
(key == 10'b0011101100) ? 46'b1010000000011001111111101010001111001011010000 :
(key == 10'b0011101101) ? 46'b1001111111000101100001001010001010111001000101 :
(key == 10'b0011101110) ? 46'b1001111101110001001011001010000110100111100011 :
(key == 10'b0011101111) ? 46'b1001111100011100111110001010000010010110101011 :
(key == 10'b0011110000) ? 46'b1001111011001000111001101001111110000110011101 :
(key == 10'b0011110001) ? 46'b1001111001110100111101101001111001110110111001 :
(key == 10'b0011110010) ? 46'b1001111000100001001001001001110101100111111101 :
(key == 10'b0011110011) ? 46'b1001110111001101011110001001110001011001101010 :
(key == 10'b0011110100) ? 46'b1001110101111001111011101001101101001011111111 :
(key == 10'b0011110101) ? 46'b1001110100100110100001001001101000111110111110 :
(key == 10'b0011110110) ? 46'b1001110011010011001111001001100100110010100101 :
(key == 10'b0011110111) ? 46'b1001110010000000000101001001100000100110110110 :
(key == 10'b0011111000) ? 46'b1001110000101101000100001001011100011011101110 :
(key == 10'b0011111001) ? 46'b1001101111011010001011101001011000010001001101 :
(key == 10'b0011111010) ? 46'b1001101110000111011011001001010100000111010110 :
(key == 10'b0011111011) ? 46'b1001101100110100110010101001001111111110000111 :
(key == 10'b0011111100) ? 46'b1001101011100010010011001001001011110101100000 :
(key == 10'b0011111101) ? 46'b1001101010001111111011001001000111101101100000 :
(key == 10'b0011111110) ? 46'b1001101000111101101011101001000011100110001000 :
(key == 10'b0011111111) ? 46'b1001100111101011100100001000111111011111010111 :
(key == 10'b0100000000) ? 46'b1001100110011001100101001000111011011001001110 :
(key == 10'b0100000001) ? 46'b1001100101000111101110101000110111010011101100 :
(key == 10'b0100000010) ? 46'b1001100011110110000000001000110011001110110010 :
(key == 10'b0100000011) ? 46'b1001100010100100011001101000101111001010011110 :
(key == 10'b0100000100) ? 46'b1001100001010010111011001000101011000110110000 :
(key == 10'b0100000101) ? 46'b1001100000000001100101001000100111000011101010 :
(key == 10'b0100000110) ? 46'b1001011110110000010111001000100011000001001011 :
(key == 10'b0100000111) ? 46'b1001011101011111010001001000011110111111010010 :
(key == 10'b0100001000) ? 46'b1001011100001110010011001000011010111101111111 :
(key == 10'b0100001001) ? 46'b1001011010111101011101001000010110111101010011 :
(key == 10'b0100001010) ? 46'b1001011001101100101111001000010010111101001101 :
(key == 10'b0100001011) ? 46'b1001011000011100001001001000001110111101101100 :
(key == 10'b0100001100) ? 46'b1001010111001011101011001000001010111110110010 :
(key == 10'b0100001101) ? 46'b1001010101111011010101001000000111000000011110 :
(key == 10'b0100001110) ? 46'b1001010100101011000111001000000011000010101111 :
(key == 10'b0100001111) ? 46'b1001010011011011000001000111111111000101100111 :
(key == 10'b0100010000) ? 46'b1001010010001011000011000111111011001001000100 :
(key == 10'b0100010001) ? 46'b1001010000111011001101000111110111001101000101 :
(key == 10'b0100010010) ? 46'b1001001111101011011110100111110011010001101100 :
(key == 10'b0100010011) ? 46'b1001001110011011110111100111101111010110111001 :
(key == 10'b0100010100) ? 46'b1001001101001100011001000111101011011100101010 :
(key == 10'b0100010101) ? 46'b1001001011111101000010000111100111100011000000 :
(key == 10'b0100010110) ? 46'b1001001010101101110011000111100011101001111011 :
(key == 10'b0100010111) ? 46'b1001001001011110101100000111011111110001011011 :
(key == 10'b0100011000) ? 46'b1001001000001111101100000111011011111001100000 :
(key == 10'b0100011001) ? 46'b1001000111000000110100100111011000000010001000 :
(key == 10'b0100011010) ? 46'b1001000101110010000100100111010100001011010100 :
(key == 10'b0100011011) ? 46'b1001000100100011011100000111010000010101000101 :
(key == 10'b0100011100) ? 46'b1001000011010100111011100111001100011111011011 :
(key == 10'b0100011101) ? 46'b1001000010000110100010100111001000101010010100 :
(key == 10'b0100011110) ? 46'b1001000000111000010001000111000100110101110001 :
(key == 10'b0100011111) ? 46'b1000111111101010000111100111000001000001110011 :
(key == 10'b0100100000) ? 46'b1000111110011100000101100110111101001110010111 :
(key == 10'b0100100001) ? 46'b1000111101001110001011000110111001011011100000 :
(key == 10'b0100100010) ? 46'b1000111100000000011000000110110101101001001100 :
(key == 10'b0100100011) ? 46'b1000111010110010101101000110110001110111011011 :
(key == 10'b0100100100) ? 46'b1000111001100101001001000110101110000110001101 :
(key == 10'b0100100101) ? 46'b1000111000010111101100100110101010010101100010 :
(key == 10'b0100100110) ? 46'b1000110111001010011000000110100110100101011010 :
(key == 10'b0100100111) ? 46'b1000110101111101001011000110100010110101110101 :
(key == 10'b0100101000) ? 46'b1000110100110000000101000110011111000110110100 :
(key == 10'b0100101001) ? 46'b1000110011100011000111000110011011011000010100 :
(key == 10'b0100101010) ? 46'b1000110010010110010000100110010111101010011000 :
(key == 10'b0100101011) ? 46'b1000110001001001100001000110010011111100111111 :
(key == 10'b0100101100) ? 46'b1000101111111100111001000110010000010000001000 :
(key == 10'b0100101101) ? 46'b1000101110110000011000100110001100100011110010 :
(key == 10'b0100101110) ? 46'b1000101101100011111111100110001000110111111111 :
(key == 10'b0100101111) ? 46'b1000101100010111101110000110000101001100101110 :
(key == 10'b0100110000) ? 46'b1000101011001011100011100110000001100001111110 :
(key == 10'b0100110001) ? 46'b1000101001111111100000100101111101110111110010 :
(key == 10'b0100110010) ? 46'b1000101000110011100100100101111010001110000110 :
(key == 10'b0100110011) ? 46'b1000100111100111110000100101110110100100111101 :
(key == 10'b0100110100) ? 46'b1000100110011100000011000101110010111100010101 :
(key == 10'b0100110101) ? 46'b1000100101010000011101000101101111010100001110 :
(key == 10'b0100110110) ? 46'b1000100100000100111110100101101011101100101000 :
(key == 10'b0100110111) ? 46'b1000100010111001100111000101101000000101100101 :
(key == 10'b0100111000) ? 46'b1000100001101110010111000101100100011111000011 :
(key == 10'b0100111001) ? 46'b1000100000100011001110000101100000111001000001 :
(key == 10'b0100111010) ? 46'b1000011111011000001100000101011101010011011111 :
(key == 10'b0100111011) ? 46'b1000011110001101010001100101011001101110100000 :
(key == 10'b0100111100) ? 46'b1000011101000010011110000101010110001010000010 :
(key == 10'b0100111101) ? 46'b1000011011110111110010000101010010100110000011 :
(key == 10'b0100111110) ? 46'b1000011010101101001100100101001111000010100101 :
(key == 10'b0100111111) ? 46'b1000011001100010101110100101001011011111101000 :
(key == 10'b0101000000) ? 46'b1000011000011000010111100101000111111101001011 :
(key == 10'b0101000001) ? 46'b1000010111001110000111100101000100011011001111 :
(key == 10'b0101000010) ? 46'b1000010110000011111110100101000000111001110010 :
(key == 10'b0101000011) ? 46'b1000010100111001111101000100111101011000110110 :
(key == 10'b0101000100) ? 46'b1000010011110000000010000100111001111000011010 :
(key == 10'b0101000101) ? 46'b1000010010100110001110100100110110011000011110 :
(key == 10'b0101000110) ? 46'b1000010001011100100010000100110010111001000001 :
(key == 10'b0101000111) ? 46'b1000010000010010111100000100101111011010000101 :
(key == 10'b0101001000) ? 46'b1000001111001001011101000100101011111011101000 :
(key == 10'b0101001001) ? 46'b1000001110000000000101100100101000011101101010 :
(key == 10'b0101001010) ? 46'b1000001100110110110100000100100101000000001100 :
(key == 10'b0101001011) ? 46'b1000001011101101101010000100100001100011001101 :
(key == 10'b0101001100) ? 46'b1000001010100100100111100100011110000110101110 :
(key == 10'b0101001101) ? 46'b1000001001011011101011000100011010101010101101 :
(key == 10'b0101001110) ? 46'b1000001000010010110101100100010111001111001100 :
(key == 10'b0101001111) ? 46'b1000000111001010000111100100010011110100001010 :
(key == 10'b0101010000) ? 46'b1000000110000001011111100100010000011001100111 :
(key == 10'b0101010001) ? 46'b1000000100111000111110100100001100111111100010 :
(key == 10'b0101010010) ? 46'b1000000011110000100101000100001001100101111101 :
(key == 10'b0101010011) ? 46'b1000000010101000010001100100000110001100110101 :
(key == 10'b0101010100) ? 46'b1000000001100000000101000100000010110100001101 :
(key == 10'b0101010101) ? 46'b1000000000010111111111100011111111011100000011 :
(key == 10'b0101010110) ? 46'b0111111111010000000000100011111100000100010111 :
(key == 10'b0101010111) ? 46'b0111111110001000001000100011111000101101001001 :
(key == 10'b0101011000) ? 46'b0111111101000000010111000011110101010110011010 :
(key == 10'b0101011001) ? 46'b0111111011111000101100100011110010000000001010 :
(key == 10'b0101011010) ? 46'b0111111010110001001000100011101110101010010110 :
(key == 10'b0101011011) ? 46'b0111111001101001101011000011101011010101000000 :
(key == 10'b0101011100) ? 46'b0111111000100010010100100011101000000000001010 :
(key == 10'b0101011101) ? 46'b0111110111011011000100100011100100101011101111 :
(key == 10'b0101011110) ? 46'b0111110110010011111011000011100001010111110011 :
(key == 10'b0101011111) ? 46'b0111110101001100111000100011011110000100010101 :
(key == 10'b0101100000) ? 46'b0111110100000101111100000011011010110001010101 :
(key == 10'b0101100001) ? 46'b0111110010111111000111000011010111011110110000 :
(key == 10'b0101100010) ? 46'b0111110001111000011000000011010100001100101010 :
(key == 10'b0101100011) ? 46'b0111110000110001101111000011010000111011000000 :
(key == 10'b0101100100) ? 46'b0111101111101011001101100011001101101001110101 :
(key == 10'b0101100101) ? 46'b0111101110100100110010000011001010011001000110 :
(key == 10'b0101100110) ? 46'b0111101101011110011101100011000111001000110100 :
(key == 10'b0101100111) ? 46'b0111101100011000001111000011000011111000111111 :
(key == 10'b0101101000) ? 46'b0111101011010010000111100011000000101001100111 :
(key == 10'b0101101001) ? 46'b0111101010001100000110000010111101011010101100 :
(key == 10'b0101101010) ? 46'b0111101001000110001011100010111010001100001101 :
(key == 10'b0101101011) ? 46'b0111101000000000010111000010110110111110001010 :
(key == 10'b0101101100) ? 46'b0111100110111010101001000010110011110000100101 :
(key == 10'b0101101101) ? 46'b0111100101110101000001100010110000100011011011 :
(key == 10'b0101101110) ? 46'b0111100100101111100000000010101101010110101110 :
(key == 10'b0101101111) ? 46'b0111100011101010000101100010101010001010011101 :
(key == 10'b0101110000) ? 46'b0111100010100100110001000010100110111110101001 :
(key == 10'b0101110001) ? 46'b0111100001011111100011100010100011110011010001 :
(key == 10'b0101110010) ? 46'b0111100000011010011011100010100000101000010100 :
(key == 10'b0101110011) ? 46'b0111011111010101011010100010011101011101110010 :
(key == 10'b0101110100) ? 46'b0111011110010000011111100010011010010011101110 :
(key == 10'b0101110101) ? 46'b0111011101001011101010100010010111001010000101 :
(key == 10'b0101110110) ? 46'b0111011100000110111100100010010100000000111000 :
(key == 10'b0101110111) ? 46'b0111011011000010010100100010010000111000000110 :
(key == 10'b0101111000) ? 46'b0111011001111101110011000010001101101111110000 :
(key == 10'b0101111001) ? 46'b0111011000111001010111000010001010100111110101 :
(key == 10'b0101111010) ? 46'b0111010111110101000010000010000111100000010110 :
(key == 10'b0101111011) ? 46'b0111010110110000110011000010000100011001010001 :
(key == 10'b0101111100) ? 46'b0111010101101100101010000010000001010010100111 :
(key == 10'b0101111101) ? 46'b0111010100101000101000000001111110001100011011 :
(key == 10'b0101111110) ? 46'b0111010011100100101011100001111011000110100111 :
(key == 10'b0101111111) ? 46'b0111010010100000110101000001111000000001010000 :
(key == 10'b0110000000) ? 46'b0111010001011101000101000001110100111100010011 :
(key == 10'b0110000001) ? 46'b0111010000011001011011100001110001110111110000 :
(key == 10'b0110000010) ? 46'b0111001111010101110111100001101110110011101001 :
(key == 10'b0110000011) ? 46'b0111001110010010011001100001101011101111111101 :
(key == 10'b0110000100) ? 46'b0111001101001111000010000001101000101100101010 :
(key == 10'b0110000101) ? 46'b0111001100001011110001000001100101101001110010 :
(key == 10'b0110000110) ? 46'b0111001011001000100101100001100010100111010110 :
(key == 10'b0110000111) ? 46'b0111001010000101100000100001011111100101010010 :
(key == 10'b0110001000) ? 46'b0111001001000010100001100001011100100011101010 :
(key == 10'b0110001001) ? 46'b0111000111111111101000000001011001100010011100 :
(key == 10'b0110001010) ? 46'b0111000110111100110101000001010110100001101000 :
(key == 10'b0110001011) ? 46'b0111000101111010001000000001010011100001001100 :
(key == 10'b0110001100) ? 46'b0111000100110111100001000001010000100001001100 :
(key == 10'b0110001101) ? 46'b0111000011110101000000000001001101100001100110 :
(key == 10'b0110001110) ? 46'b0111000010110010100101000001001010100010011010 :
(key == 10'b0110001111) ? 46'b0111000001110000010000000001000111100011101000 :
(key == 10'b0110010000) ? 46'b0111000000101110000000100001000100100101010000 :
(key == 10'b0110010001) ? 46'b0110111111101011110111100001000001100111001111 :
(key == 10'b0110010010) ? 46'b0110111110101001110100000000111110101001101011 :
(key == 10'b0110010011) ? 46'b0110111101100111110111000000111011101100011110 :
(key == 10'b0110010100) ? 46'b0110111100100110000000000000111000101111101011 :
(key == 10'b0110010101) ? 46'b0110111011100100001110000000110101110011010010 :
(key == 10'b0110010110) ? 46'b0110111010100010100010100000110010110111010010 :
(key == 10'b0110010111) ? 46'b0110111001100000111100100000101111111011101011 :
(key == 10'b0110011000) ? 46'b0110111000011111011101000000101101000000011101 :
(key == 10'b0110011001) ? 46'b0110110111011110000011000000101010000101101000 :
(key == 10'b0110011010) ? 46'b0110110110011100101110100000100111001011001101 :
(key == 10'b0110011011) ? 46'b0110110101011011100000100000100100010001001010 :
(key == 10'b0110011100) ? 46'b0110110100011010011000000000100001010111011111 :
(key == 10'b0110011101) ? 46'b0110110011011001010101000000011110011110001111 :
(key == 10'b0110011110) ? 46'b0110110010011000011000000000011011100101010111 :
(key == 10'b0110011111) ? 46'b0110110001010111100001000000011000101100110111 :
(key == 10'b0110100000) ? 46'b0110110000010110101111100000010101110100101111 :
(key == 10'b0110100001) ? 46'b0110101111010110000100000000010010111101000010 :
(key == 10'b0110100010) ? 46'b0110101110010101011110000000010000000101101010 :
(key == 10'b0110100011) ? 46'b0110101101010100111110000000001101001110101101 :
(key == 10'b0110100100) ? 46'b0110101100010100100011100000001010011000001000 :
(key == 10'b0110100101) ? 46'b0110101011010100001110100000000111100001111010 :
(key == 10'b0110100110) ? 46'b0110101010010011111111100000000100101100000100 :
(key == 10'b0110100111) ? 46'b0110101001010011110110100000000001110110101000 :
(key == 10'b0110101000) ? 46'b0110101000010011110010111111111110000011000100 :
(key == 10'b0110101001) ? 46'b0110100111010011110100111111111000011001101100 :
(key == 10'b0110101010) ? 46'b0110100110010011111100011111110010110001000010 :
(key == 10'b0110101011) ? 46'b0110100101010100001001111111101101001001000111 :
(key == 10'b0110101100) ? 46'b0110100100010100011100111111100111100001111100 :
(key == 10'b0110101101) ? 46'b0110100011010100110100111111100001111011100001 :
(key == 10'b0110101110) ? 46'b0110100010010101010011011111011100010101110110 :
(key == 10'b0110101111) ? 46'b0110100001010101110110111111010110110000110110 :
(key == 10'b0110110000) ? 46'b0110100000010110011111111111010001001100101011 :
(key == 10'b0110110001) ? 46'b0110011111010111001110111111001011101001001100 :
(key == 10'b0110110010) ? 46'b0110011110011000000010111111000110000110011011 :
(key == 10'b0110110011) ? 46'b0110011101011000111100111111000000100100011000 :
(key == 10'b0110110100) ? 46'b0110011100011001111100011110111011000011000111 :
(key == 10'b0110110101) ? 46'b0110011011011011000001011110110101100010100001 :
(key == 10'b0110110110) ? 46'b0110011010011100001011111110110000000010101001 :
(key == 10'b0110110111) ? 46'b0110011001011101011011111110101010100011100011 :
(key == 10'b0110111000) ? 46'b0110011000011110110001011110100101000101000111 :
(key == 10'b0110111001) ? 46'b0110010111100000001011111110011111100111011101 :
(key == 10'b0110111010) ? 46'b0110010110100001101100111110011010001010011110 :
(key == 10'b0110111011) ? 46'b0110010101100011010010011110010100101110001100 :
(key == 10'b0110111100) ? 46'b0110010100100100111101111110001111010010101001 :
(key == 10'b0110111101) ? 46'b0110010011100110101110011110001001110111110011 :
(key == 10'b0110111110) ? 46'b0110010010101000100100011110000100011101101001 :
(key == 10'b0110111111) ? 46'b0110010001101010100000011101111111000100001111 :
(key == 10'b0111000000) ? 46'b0110010000101100100000111101111001101011011111 :
(key == 10'b0111000001) ? 46'b0110001111101110100111011101110100010011011110 :
(key == 10'b0111000010) ? 46'b0110001110110000110010111101101110111100001001 :
(key == 10'b0111000011) ? 46'b0110001101110011000100011101101001100101100000 :
(key == 10'b0111000100) ? 46'b0110001100110101011010111101100100001111100110 :
(key == 10'b0111000101) ? 46'b0110001011110111110110011101011110111010010101 :
(key == 10'b0111000110) ? 46'b0110001010111010010111011101011001100101110011 :
(key == 10'b0111000111) ? 46'b0110001001111100111101111101010100010001111100 :
(key == 10'b0111001000) ? 46'b0110001000111111101001111101001110111110110010 :
(key == 10'b0111001001) ? 46'b0110001000000010011010011101001001101100010010 :
(key == 10'b0111001010) ? 46'b0110000111000101010000111101000100011010100000 :
(key == 10'b0111001011) ? 46'b0110000110001000001100011100111111001001010111 :
(key == 10'b0111001100) ? 46'b0110000101001011001101011100111001111000111011 :
(key == 10'b0111001101) ? 46'b0110000100001110010011011100110100101001001101 :
(key == 10'b0111001110) ? 46'b0110000011010001011110111100101111011010001000 :
(key == 10'b0111001111) ? 46'b0110000010010100101111011100101010001011101101 :
(key == 10'b0111010000) ? 46'b0110000001011000000101011100100100111101111111 :
(key == 10'b0111010001) ? 46'b0110000000011011100000011100011111110000111011 :
(key == 10'b0111010010) ? 46'b0101111111011111000000011100011010100100100011 :
(key == 10'b0111010011) ? 46'b0101111110100010100101111100010101011000110101 :
(key == 10'b0111010100) ? 46'b0101111101100110010000011100010000001101110001 :
(key == 10'b0111010101) ? 46'b0101111100101010000000011100001011000011011001 :
(key == 10'b0111010110) ? 46'b0101111011101101110101011100000101111001101011 :
(key == 10'b0111010111) ? 46'b0101111010110001101111011100000000110000101000 :
(key == 10'b0111011000) ? 46'b0101111001110101101110111011111011101000001101 :
(key == 10'b0111011001) ? 46'b0101111000111001110010111011110110100000011110 :
(key == 10'b0111011010) ? 46'b0101110111111101111100011011110001011001011000 :
(key == 10'b0111011011) ? 46'b0101110111000010001010111011101100010010111011 :
(key == 10'b0111011100) ? 46'b0101110110000110011110111011100111001101001011 :
(key == 10'b0111011101) ? 46'b0101110101001010110111011011100010001000000011 :
(key == 10'b0111011110) ? 46'b0101110100001111010101011011011101000011100010 :
(key == 10'b0111011111) ? 46'b0101110011010011111000011011010111111111101101 :
(key == 10'b0111100000) ? 46'b0101110010011000100000011011010010111100100001 :
(key == 10'b0111100001) ? 46'b0101110001011101001101011011001101111010000000 :
(key == 10'b0111100010) ? 46'b0101110000100001111111011011001000111000000110 :
(key == 10'b0111100011) ? 46'b0101101111100110110110111011000011110110110100 :
(key == 10'b0111100100) ? 46'b0101101110101011110010111010111110110110001011 :
(key == 10'b0111100101) ? 46'b0101101101110000110011111010111001110110001110 :
(key == 10'b0111100110) ? 46'b0101101100110101111010011010110100110110110111 :
(key == 10'b0111100111) ? 46'b0101101011111011000101011010101111111000001000 :
(key == 10'b0111101000) ? 46'b0101101011000000010101011010101010111010000010 :
(key == 10'b0111101001) ? 46'b0101101010000101101010011010100101111100100111 :
(key == 10'b0111101010) ? 46'b0101101001001011000100111010100000111111110010 :
(key == 10'b0111101011) ? 46'b0101101000010000100011111010011100000011100101 :
(key == 10'b0111101100) ? 46'b0101100111010110000111011010010111000111111110 :
(key == 10'b0111101101) ? 46'b0101100110011011110000011010010010001101000010 :
(key == 10'b0111101110) ? 46'b0101100101100001011110011010001101010010101111 :
(key == 10'b0111101111) ? 46'b0101100100100111010000111010001000011001000000 :
(key == 10'b0111110000) ? 46'b0101100011101101001000011010000011011111111010 :
(key == 10'b0111110001) ? 46'b0101100010110011000100111001111110100111011100 :
(key == 10'b0111110010) ? 46'b0101100001111001000110011001111001101111100110 :
(key == 10'b0111110011) ? 46'b0101100000111111001100011001110100111000010110 :
(key == 10'b0111110100) ? 46'b0101100000000101010111111001110000000001101101 :
(key == 10'b0111110101) ? 46'b0101011111001011100111111001101011001011101100 :
(key == 10'b0111110110) ? 46'b0101011110010001111100011001100110010110010001 :
(key == 10'b0111110111) ? 46'b0101011101011000010110011001100001100001011101 :
(key == 10'b0111111000) ? 46'b0101011100011110110100111001011100101101010001 :
(key == 10'b0111111001) ? 46'b0101011011100101010111111001010111111001101100 :
(key == 10'b0111111010) ? 46'b0101011010101100000000011001010011000110101101 :
(key == 10'b0111111011) ? 46'b0101011001110010101100111001001110010100010011 :
(key == 10'b0111111100) ? 46'b0101011000111001011110011001001001100010100000 :
(key == 10'b0111111101) ? 46'b0101011000000000010100111001000100110001010100 :
(key == 10'b0111111110) ? 46'b0101010111000111010000011001000000000000101101 :
(key == 10'b0111111111) ? 46'b0101010110001110010000011000111011010000101110 :
(key == 10'b1000000000) ? 46'b0101010101010101010100111000110110100001010011 :
(key == 10'b1000000001) ? 46'b0101010100011100011110011000110001110010100000 :
(key == 10'b1000000010) ? 46'b0101010011100011101100111000101101000100010001 :
(key == 10'b1000000011) ? 46'b0101010010101010111111011000101000010110101010 :
(key == 10'b1000000100) ? 46'b0101010001110010010111011000100011101001100110 :
(key == 10'b1000000101) ? 46'b0101010000111001110011111000011110111101001000 :
(key == 10'b1000000110) ? 46'b0101010000000001010100111000011010010001010000 :
(key == 10'b1000000111) ? 46'b0101001111001000111010011000010101100101111101 :
(key == 10'b1000001000) ? 46'b0101001110010000100100111000010000111011001101 :
(key == 10'b1000001001) ? 46'b0101001101011000010011111000001100010001000101 :
(key == 10'b1000001010) ? 46'b0101001100100000000111111000000111100111100001 :
(key == 10'b1000001011) ? 46'b0101001011101000000000011000000010111110100100 :
(key == 10'b1000001100) ? 46'b0101001010101111111101010111111110010110001000 :
(key == 10'b1000001101) ? 46'b0101001001110111111110110111111001101110010011 :
(key == 10'b1000001110) ? 46'b0101001001000000000100110111110101000111000010 :
(key == 10'b1000001111) ? 46'b0101001000001000001111110111110000100000011000 :
(key == 10'b1000010000) ? 46'b0101000111010000011111010111101011111010001110 :
(key == 10'b1000010001) ? 46'b0101000110011000110011010111100111010100101100 :
(key == 10'b1000010010) ? 46'b0101000101100001001100010111100010101111101101 :
(key == 10'b1000010011) ? 46'b0101000100101001101001010111011110001011010001 :
(key == 10'b1000010100) ? 46'b0101000011110010001011010111011001100111011010 :
(key == 10'b1000010101) ? 46'b0101000010111010110001110111010101000100001001 :
(key == 10'b1000010110) ? 46'b0101000010000011011100110111010000100001011001 :
(key == 10'b1000010111) ? 46'b0101000001001100001100010111001011111111001111 :
(key == 10'b1000011000) ? 46'b0101000000010100111111110111000111011101100110 :
(key == 10'b1000011001) ? 46'b0100111111011101111000110111000010111100100011 :
(key == 10'b1000011010) ? 46'b0100111110100110110101110110111110011100000001 :
(key == 10'b1000011011) ? 46'b0100111101101111110111010110111001111100000101 :
(key == 10'b1000011100) ? 46'b0100111100111000111101010110110101011100101100 :
(key == 10'b1000011101) ? 46'b0100111100000010000111110110110000111101110100 :
(key == 10'b1000011110) ? 46'b0100111011001011010110110110101100011111100010 :
(key == 10'b1000011111) ? 46'b0100111010010100101010010110101000000001110000 :
(key == 10'b1000100000) ? 46'b0100111001011110000010010110100011100100100100 :
(key == 10'b1000100001) ? 46'b0100111000100111011110110110011111000111111001 :
(key == 10'b1000100010) ? 46'b0100110111110000111111110110011010101011110001 :
(key == 10'b1000100011) ? 46'b0100110110111010100101010110010110010000001100 :
(key == 10'b1000100100) ? 46'b0100110110000100001110110110010001110101001010 :
(key == 10'b1000100101) ? 46'b0100110101001101111100110110001101011010101011 :
(key == 10'b1000100110) ? 46'b0100110100010111101111010110001001000000101100 :
(key == 10'b1000100111) ? 46'b0100110011100001100110010110000100100111010010 :
(key == 10'b1000101000) ? 46'b0100110010101011100001110110000000001110011001 :
(key == 10'b1000101001) ? 46'b0100110001110101100001110101111011110110000011 :
(key == 10'b1000101010) ? 46'b0100110000111111100101110101110111011110001111 :
(key == 10'b1000101011) ? 46'b0100110000001001101110010101110011000110111100 :
(key == 10'b1000101100) ? 46'b0100101111010011111011010101101110110000001011 :
(key == 10'b1000101101) ? 46'b0100101110011110001100110101101010011001111100 :
(key == 10'b1000101110) ? 46'b0100101101101000100001110101100110000100010000 :
(key == 10'b1000101111) ? 46'b0100101100110010111011110101100001101111000101 :
(key == 10'b1000110000) ? 46'b0100101011111101011010010101011101011010011011 :
(key == 10'b1000110001) ? 46'b0100101011000111111100110101011001000110010010 :
(key == 10'b1000110010) ? 46'b0100101010010010100011110101010100110010101011 :
(key == 10'b1000110011) ? 46'b0100101001011101001110110101010000011111100110 :
(key == 10'b1000110100) ? 46'b0100101000100111111110110101001100001101000001 :
(key == 10'b1000110101) ? 46'b0100100111110010110010010101000111111010111110 :
(key == 10'b1000110110) ? 46'b0100100110111101101010010101000011101001011101 :
(key == 10'b1000110111) ? 46'b0100100110001000100110110100111111011000011010 :
(key == 10'b1000111000) ? 46'b0100100101010011100111010100111011000111111011 :
(key == 10'b1000111001) ? 46'b0100100100011110101100010100110110110111111011 :
(key == 10'b1000111010) ? 46'b0100100011101001110101010100110010101000011100 :
(key == 10'b1000111011) ? 46'b0100100010110101000010110100101110011001011110 :
(key == 10'b1000111100) ? 46'b0100100010000000010100010100101010001011000010 :
(key == 10'b1000111101) ? 46'b0100100001001011101010010100100101111101000101 :
(key == 10'b1000111110) ? 46'b0100100000010111000100010100100001101111101000 :
(key == 10'b1000111111) ? 46'b0100011111100010100010110100011101100010101101 :
(key == 10'b1001000000) ? 46'b0100011110101110000100110100011001010110010000 :
(key == 10'b1001000001) ? 46'b0100011101111001101011110100010101001010010011 :
(key == 10'b1001000010) ? 46'b0100011101000101010110010100010000111110111000 :
(key == 10'b1001000011) ? 46'b0100011100010001000101110100001100110011111100 :
(key == 10'b1001000100) ? 46'b0100011011011100111000110100001000101001100010 :
(key == 10'b1001000101) ? 46'b0100011010101000101111110100000100011111100110 :
(key == 10'b1001000110) ? 46'b0100011001110100101011010100000000010110001010 :
(key == 10'b1001000111) ? 46'b0100011001000000101011010011111100001101001100 :
(key == 10'b1001001000) ? 46'b0100011000001100101110110011111000000100110000 :
(key == 10'b1001001001) ? 46'b0100010111011000110110110011110011111100110011 :
(key == 10'b1001001010) ? 46'b0100010110100101000010110011101111110101010101 :
(key == 10'b1001001011) ? 46'b0100010101110001010011010011101011101110011000 :
(key == 10'b1001001100) ? 46'b0100010100111101100111010011100111100111110111 :
(key == 10'b1001001101) ? 46'b0100010100001001111111110011100011100001111000 :
(key == 10'b1001001110) ? 46'b0100010011010110011100010011011111011100010111 :
(key == 10'b1001001111) ? 46'b0100010010100010111100110011011011010111010111 :
(key == 10'b1001010000) ? 46'b0100010001101111100001010011010111010010110100 :
(key == 10'b1001010001) ? 46'b0100010000111100001001110011010011001110101111 :
(key == 10'b1001010010) ? 46'b0100010000001000110110110011001111001011001011 :
(key == 10'b1001010011) ? 46'b0100001111010101100111110011001011001000000110 :
(key == 10'b1001010100) ? 46'b0100001110100010011100110011000111000101011100 :
(key == 10'b1001010101) ? 46'b0100001101101111010101010011000011000011010100 :
(key == 10'b1001010110) ? 46'b0100001100111100010010010010111111000001101010 :
(key == 10'b1001010111) ? 46'b0100001100001001010011010010111011000000011110 :
(key == 10'b1001011000) ? 46'b0100001011010110011000010010110110111111110001 :
(key == 10'b1001011001) ? 46'b0100001010100011100001010010110010111111100010 :
(key == 10'b1001011010) ? 46'b0100001001110000101110010010101110111111110001 :
(key == 10'b1001011011) ? 46'b0100001000111101111111010010101011000000011110 :
(key == 10'b1001011100) ? 46'b0100001000001011010100010010100111000001101001 :
(key == 10'b1001011101) ? 46'b0100000111011000101101010010100011000011010011 :
(key == 10'b1001011110) ? 46'b0100000110100110001010010010011111000101011011 :
(key == 10'b1001011111) ? 46'b0100000101110011101011010010011011001000000000 :
(key == 10'b1001100000) ? 46'b0100000101000001010000010010010111001011000010 :
(key == 10'b1001100001) ? 46'b0100000100001110111000110010010011001110100011 :
(key == 10'b1001100010) ? 46'b0100000011011100100101110010001111010010100011 :
(key == 10'b1001100011) ? 46'b0100000010101010010110010010001011010110111110 :
(key == 10'b1001100100) ? 46'b0100000001111000001011010010000111011011110111 :
(key == 10'b1001100101) ? 46'b0100000001000110000011010010000011100001001110 :
(key == 10'b1001100110) ? 46'b0100000000010100000000010001111111100111000011 :
(key == 10'b1001100111) ? 46'b0011111111100010000000110001111011101101010101 :
(key == 10'b1001101000) ? 46'b0011111110110000000100110001110111110100000010 :
(key == 10'b1001101001) ? 46'b0011111101111110001100110001110011111011001110 :
(key == 10'b1001101010) ? 46'b0011111101001100011000110001110000000010110111 :
(key == 10'b1001101011) ? 46'b0011111100011010101000110001101100001010111101 :
(key == 10'b1001101100) ? 46'b0011111011101000111100110001101000010011100001 :
(key == 10'b1001101101) ? 46'b0011111010110111010100010001100100011100100001 :
(key == 10'b1001101110) ? 46'b0011111010000101101111110001100000100101111101 :
(key == 10'b1001101111) ? 46'b0011111001010100001111110001011100101111110111 :
(key == 10'b1001110000) ? 46'b0011111000100010110010110001011000111010001100 :
(key == 10'b1001110001) ? 46'b0011110111110001011001110001010101000100111111 :
(key == 10'b1001110010) ? 46'b0011110111000000000100110001010001010000001111 :
(key == 10'b1001110011) ? 46'b0011110110001110110011110001001101011011111010 :
(key == 10'b1001110100) ? 46'b0011110101011101100110010001001001101000000010 :
(key == 10'b1001110101) ? 46'b0011110100101100011100010001000101110100100101 :
(key == 10'b1001110110) ? 46'b0011110011111011010110110001000010000001100111 :
(key == 10'b1001110111) ? 46'b0011110011001010010100110000111110001111000010 :
(key == 10'b1001111000) ? 46'b0011110010011001010110010000111010011100111100 :
(key == 10'b1001111001) ? 46'b0011110001101000011011110000110110101011010001 :
(key == 10'b1001111010) ? 46'b0011110000110111100101010000110010111010000001 :
(key == 10'b1001111011) ? 46'b0011110000000110110010010000101111001001001110 :
(key == 10'b1001111100) ? 46'b0011101111010110000011010000101011011000110101 :
(key == 10'b1001111101) ? 46'b0011101110100101010111110000100111101000111010 :
(key == 10'b1001111110) ? 46'b0011101101110100110000010000100011111001011011 :
(key == 10'b1001111111) ? 46'b0011101101000100001100010000100000001010010111 :
(key == 10'b1010000000) ? 46'b0011101100010011101011110000011100011011101101 :
(key == 10'b1010000001) ? 46'b0011101011100011001111110000011000101101100000 :
(key == 10'b1010000010) ? 46'b0011101010110010110111010000010100111111101101 :
(key == 10'b1010000011) ? 46'b0011101010000010100001110000010001010010010111 :
(key == 10'b1010000100) ? 46'b0011101001010010010000110000001101100101011100 :
(key == 10'b1010000101) ? 46'b0011101000100010000011010000001001111000111101 :
(key == 10'b1010000110) ? 46'b0011100111110001111001010000000110001100111000 :
(key == 10'b1010000111) ? 46'b0011100111000001110011010000000010100001001110 :
(key == 10'b1010001000) ? 46'b0011100110010001110000001111111110110110000000 :
(key == 10'b1010001001) ? 46'b0011100101100001110001101111111011001011001100 :
(key == 10'b1010001010) ? 46'b0011100100110001110110101111110111100000110011 :
(key == 10'b1010001011) ? 46'b0011100100000001111110101111110011110110110011 :
(key == 10'b1010001100) ? 46'b0011100011010010001011001111110000001101010000 :
(key == 10'b1010001101) ? 46'b0011100010100010011011001111101100100100001010 :
(key == 10'b1010001110) ? 46'b0011100001110010101110001111101000111011011011 :
(key == 10'b1010001111) ? 46'b0011100001000011000101001111100101010011001000 :
(key == 10'b1010010000) ? 46'b0011100000010011100000001111100001101011010000 :
(key == 10'b1010010001) ? 46'b0011011111100011111110101111011110000011110001 :
(key == 10'b1010010010) ? 46'b0011011110110100100000001111011010011100101110 :
(key == 10'b1010010011) ? 46'b0011011110000101000101101111010110110110000011 :
(key == 10'b1010010100) ? 46'b0011011101010101101111001111010011001111110100 :
(key == 10'b1010010101) ? 46'b0011011100100110011011101111001111101001111111 :
(key == 10'b1010010110) ? 46'b0011011011110111001100001111001100000100100110 :
(key == 10'b1010010111) ? 46'b0011011011001000000000001111001000011111100100 :
(key == 10'b1010011000) ? 46'b0011011010011000110111101111000100111010111111 :
(key == 10'b1010011001) ? 46'b0011011001101001110010101111000001010110110000 :
(key == 10'b1010011010) ? 46'b0011011000111010110001001110111101110010111110 :
(key == 10'b1010011011) ? 46'b0011011000001011110011001110111010001111100101 :
(key == 10'b1010011100) ? 46'b0011010111011100111001001110110110101100100110 :
(key == 10'b1010011101) ? 46'b0011010110101110000010101110110011001010000000 :
(key == 10'b1010011110) ? 46'b0011010101111111001111001110101111100111110110 :
(key == 10'b1010011111) ? 46'b0011010101010000011111101110101100000110000100 :
(key == 10'b1010100000) ? 46'b0011010100100001110011101110101000100100101010 :
(key == 10'b1010100001) ? 46'b0011010011110011001011001110100101000011101101 :
(key == 10'b1010100010) ? 46'b0011010011000100100101101110100001100011000110 :
(key == 10'b1010100011) ? 46'b0011010010010110000100001110011110000010111001 :
(key == 10'b1010100100) ? 46'b0011010001100111100110001110011010100011000111 :
(key == 10'b1010100101) ? 46'b0011010000111001001011101110010111000011101101 :
(key == 10'b1010100110) ? 46'b0011010000001010110100101110010011100100101110 :
(key == 10'b1010100111) ? 46'b0011001111011100100001001110010000000110000101 :
(key == 10'b1010101000) ? 46'b0011001110101110010001001110001100100111110110 :
(key == 10'b1010101001) ? 46'b0011001110000000000100101110001001001010000001 :
(key == 10'b1010101010) ? 46'b0011001101010001111011101110000101101100100110 :
(key == 10'b1010101011) ? 46'b0011001100100011110101101110000010001111100011 :
(key == 10'b1010101100) ? 46'b0011001011110101110011101101111110110010111000 :
(key == 10'b1010101101) ? 46'b0011001011000111110100101101111011010110100100 :
(key == 10'b1010101110) ? 46'b0011001010011001111001001101110111111010101100 :
(key == 10'b1010101111) ? 46'b0011001001101100000001101101110100011111001100 :
(key == 10'b1010110000) ? 46'b0011001000111110001100101101110001000100000011 :
(key == 10'b1010110001) ? 46'b0011001000010000011011101101101101101001010101 :
(key == 10'b1010110010) ? 46'b0011000111100010101110001101101010001110111110 :
(key == 10'b1010110011) ? 46'b0011000110110101000100001101100110110101000000 :
(key == 10'b1010110100) ? 46'b0011000110000111011101001101100011011011011000 :
(key == 10'b1010110101) ? 46'b0011000101011001111001101101100000000010001011 :
(key == 10'b1010110110) ? 46'b0011000100101100011001101101011100101001010101 :
(key == 10'b1010110111) ? 46'b0011000011111110111101001101011001010000111000 :
(key == 10'b1010111000) ? 46'b0011000011010001100011101101010101111000110011 :
(key == 10'b1010111001) ? 46'b0011000010100100001101101101010010100001000111 :
(key == 10'b1010111010) ? 46'b0011000001110110111011101101001111001001110001 :
(key == 10'b1010111011) ? 46'b0011000001001001101100001101001011110010110100 :
(key == 10'b1010111100) ? 46'b0011000000011100100000101101001000011100001111 :
(key == 10'b1010111101) ? 46'b0010111111101111011000001101000101000110000001 :
(key == 10'b1010111110) ? 46'b0010111111000010010011001101000001110000001110 :
(key == 10'b1010111111) ? 46'b0010111110010101010001001100111110011010101110 :
(key == 10'b1011000000) ? 46'b0010111101101000010010101100111011000101101001 :
(key == 10'b1011000001) ? 46'b0010111100111011010111101100110111110000111011 :
(key == 10'b1011000010) ? 46'b0010111100001110100000001100110100011100100101 :
(key == 10'b1011000011) ? 46'b0010111011100001101011101100110001001000100100 :
(key == 10'b1011000100) ? 46'b0010111010110100111010001100101101110100111101 :
(key == 10'b1011000101) ? 46'b0010111010001000001100101100101010100001101101 :
(key == 10'b1011000110) ? 46'b0010111001011011100001101100100111001110110100 :
(key == 10'b1011000111) ? 46'b0010111000101110111010101100100011111100010011 :
(key == 10'b1011001000) ? 46'b0010111000000010010110101100100000101010000111 :
(key == 10'b1011001001) ? 46'b0010110111010101110110001100011101011000010100 :
(key == 10'b1011001010) ? 46'b0010110110101001011000101100011010000110111010 :
(key == 10'b1011001011) ? 46'b0010110101111100111110101100010110110101110101 :
(key == 10'b1011001100) ? 46'b0010110101010000100111101100010011100101000110 :
(key == 10'b1011001101) ? 46'b0010110100100100010100001100010000010100110001 :
(key == 10'b1011001110) ? 46'b0010110011111000000011101100001101000100110000 :
(key == 10'b1011001111) ? 46'b0010110011001011110110101100001001110101000111 :
(key == 10'b1011010000) ? 46'b0010110010011111101101001100000110100101110110 :
(key == 10'b1011010001) ? 46'b0010110001110011100110001100000011010110111011 :
(key == 10'b1011010010) ? 46'b0010110001000111100010101100000000001000010101 :
(key == 10'b1011010011) ? 46'b0010110000011011100011001011111100111010000111 :
(key == 10'b1011010100) ? 46'b0010101111101111100110001011111001101100010001 :
(key == 10'b1011010101) ? 46'b0010101111000011101100001011110110011110110001 :
(key == 10'b1011010110) ? 46'b0010101110010111110101101011110011010001100111 :
(key == 10'b1011010111) ? 46'b0010101101101100000010101011110000000100110010 :
(key == 10'b1011011000) ? 46'b0010101101000000010010001011101100111000010111 :
(key == 10'b1011011001) ? 46'b0010101100010100100101101011101001101100001111 :
(key == 10'b1011011010) ? 46'b0010101011101000111011101011100110100000011111 :
(key == 10'b1011011011) ? 46'b0010101010111101010101001011100011010101000100 :
(key == 10'b1011011100) ? 46'b0010101010010001110010001011100000001001111111 :
(key == 10'b1011011101) ? 46'b0010101001100110010001101011011100111111010010 :
(key == 10'b1011011110) ? 46'b0010101000111010110101001011011001110100111010 :
(key == 10'b1011011111) ? 46'b0010101000001111011011001011010110101010111010 :
(key == 10'b1011100000) ? 46'b0010100111100100000100001011010011100001001111 :
(key == 10'b1011100001) ? 46'b0010100110111000110001001011010000010111111001 :
(key == 10'b1011100010) ? 46'b0010100110001101100000101011001101001110111000 :
(key == 10'b1011100011) ? 46'b0010100101100010010011001011001010000110001111 :
(key == 10'b1011100100) ? 46'b0010100100110111001001001011000110111101111100 :
(key == 10'b1011100101) ? 46'b0010100100001100000010001011000011110101111101 :
(key == 10'b1011100110) ? 46'b0010100011100000111110101011000000101110010110 :
(key == 10'b1011100111) ? 46'b0010100010110101111101101010111101100111000010 :
(key == 10'b1011101000) ? 46'b0010100010001011000000001010111010100000000101 :
(key == 10'b1011101001) ? 46'b0010100001100000000101101010110111011001011101 :
(key == 10'b1011101010) ? 46'b0010100000110101001110001010110100010011001010 :
(key == 10'b1011101011) ? 46'b0010100000001010011001101010110001001101001111 :
(key == 10'b1011101100) ? 46'b0010011111011111101000101010101110000111101001 :
(key == 10'b1011101101) ? 46'b0010011110110100111010001010101011000010010101 :
(key == 10'b1011101110) ? 46'b0010011110001010001111101010100111111101011001 :
(key == 10'b1011101111) ? 46'b0010011101011111100111101010100100111000110100 :
(key == 10'b1011110000) ? 46'b0010011100110101000010101010100001110100100001 :
(key == 10'b1011110001) ? 46'b0010011100001010100001001010011110110000100100 :
(key == 10'b1011110010) ? 46'b0010011011100000000010001010011011101100111110 :
(key == 10'b1011110011) ? 46'b0010011010110101100110001010011000101001101100 :
(key == 10'b1011110100) ? 46'b0010011010001011001101101010010101100110101101 :
(key == 10'b1011110101) ? 46'b0010011001100000111000001010010010100100000101 :
(key == 10'b1011110110) ? 46'b0010011000110110100101101010001111100001110010 :
(key == 10'b1011110111) ? 46'b0010011000001100010110001010001100011111110100 :
(key == 10'b1011111000) ? 46'b0010010111100010001001101010001001011110001010 :
(key == 10'b1011111001) ? 46'b0010010110111000000000001010000110011100110101 :
(key == 10'b1011111010) ? 46'b0010010110001101111001101010000011011011110101 :
(key == 10'b1011111011) ? 46'b0010010101100011110110001010000000011011001001 :
(key == 10'b1011111100) ? 46'b0010010100111001110101101001111101011010110101 :
(key == 10'b1011111101) ? 46'b0010010100001111111000001001111010011010110010 :
(key == 10'b1011111110) ? 46'b0010010011100101111110001001110111011011000101 :
(key == 10'b1011111111) ? 46'b0010010010111100000110101001110100011011101100 :
(key == 10'b1100000000) ? 46'b0010010010010010010010001001110001011100100111 :
(key == 10'b1100000001) ? 46'b0010010001101000100000101001101110011101110111 :
(key == 10'b1100000010) ? 46'b0010010000111110110010001001101011011111011011 :
(key == 10'b1100000011) ? 46'b0010010000010101000110101001101000100001010100 :
(key == 10'b1100000100) ? 46'b0010001111101011011110001001100101100011100010 :
(key == 10'b1100000101) ? 46'b0010001111000001111000101001100010100110000100 :
(key == 10'b1100000110) ? 46'b0010001110011000010110001001011111101000111010 :
(key == 10'b1100000111) ? 46'b0010001101101110110110001001011100101100000010 :
(key == 10'b1100001000) ? 46'b0010001101000101011001101001011001101111100001 :
(key == 10'b1100001001) ? 46'b0010001100011100000000001001010110110011010010 :
(key == 10'b1100001010) ? 46'b0010001011110010101001001001010011110111011010 :
(key == 10'b1100001011) ? 46'b0010001011001001010101001001010000111011110100 :
(key == 10'b1100001100) ? 46'b0010001010100000000100101001001110000000100010 :
(key == 10'b1100001101) ? 46'b0010001001110110110110001001001011000101100100 :
(key == 10'b1100001110) ? 46'b0010001001001101101011001001001000001010111010 :
(key == 10'b1100001111) ? 46'b0010001000100100100011001001000101010000100011 :
(key == 10'b1100010000) ? 46'b0010000111111011011110001001000010010110100010 :
(key == 10'b1100010001) ? 46'b0010000111010010011011001000111111011100110010 :
(key == 10'b1100010010) ? 46'b0010000110101001011100001000111100100011010111 :
(key == 10'b1100010011) ? 46'b0010000110000000011111101000111001101010010000 :
(key == 10'b1100010100) ? 46'b0010000101010111100101101000110110110001011011 :
(key == 10'b1100010101) ? 46'b0010000100101110101111001000110011111000111100 :
(key == 10'b1100010110) ? 46'b0010000100000101111011001000110001000000101111 :
(key == 10'b1100010111) ? 46'b0010000011011101001010001000101110001000110111 :
(key == 10'b1100011000) ? 46'b0010000010110100011100001000101011010001001111 :
(key == 10'b1100011001) ? 46'b0010000010001011110000101000101000011001111100 :
(key == 10'b1100011010) ? 46'b0010000001100011001000101000100101100010111101 :
(key == 10'b1100011011) ? 46'b0010000000111010100010101000100010101100010010 :
(key == 10'b1100011100) ? 46'b0010000000010010000000001000011111110101111010 :
(key == 10'b1100011101) ? 46'b0001111111101001100000001000011100111111110101 :
(key == 10'b1100011110) ? 46'b0001111111000001000011001000011010001010000011 :
(key == 10'b1100011111) ? 46'b0001111110011000101001001000010111010100100011 :
(key == 10'b1100100000) ? 46'b0001111101110000010001101000010100011111010110 :
(key == 10'b1100100001) ? 46'b0001111101000111111101001000010001101010011110 :
(key == 10'b1100100010) ? 46'b0001111100011111101011101000001110110101111001 :
(key == 10'b1100100011) ? 46'b0001111011110111011100101000001100000001100110 :
(key == 10'b1100100100) ? 46'b0001111011001111010000101000001001001101100110 :
(key == 10'b1100100101) ? 46'b0001111010100111000111101000000110011001111000 :
(key == 10'b1100100110) ? 46'b0001111001111111000001001000000011100110011110 :
(key == 10'b1100100111) ? 46'b0001111001010110111101101000000000110011011000 :
(key == 10'b1100101000) ? 46'b0001111000101110111100100111111110000000100010 :
(key == 10'b1100101001) ? 46'b0001111000000110111110100111111011001110000001 :
(key == 10'b1100101010) ? 46'b0001110111011111000011000111111000011011110001 :
(key == 10'b1100101011) ? 46'b0001110110110111001011000111110101101001110101 :
(key == 10'b1100101100) ? 46'b0001110110001111010101000111110010111000001001 :
(key == 10'b1100101101) ? 46'b0001110101100111100010100111110000000110110010 :
(key == 10'b1100101110) ? 46'b0001110100111111110010000111101101010101101110 :
(key == 10'b1100101111) ? 46'b0001110100011000000101000111101010100100111011 :
(key == 10'b1100110000) ? 46'b0001110011110000011010100111100111110100011100 :
(key == 10'b1100110001) ? 46'b0001110011001000110010100111100101000100001110 :
(key == 10'b1100110010) ? 46'b0001110010100001001101100111100010010100010010 :
(key == 10'b1100110011) ? 46'b0001110001111001101011000111011111100100101000 :
(key == 10'b1100110100) ? 46'b0001110001010010001011100111011100110101010011 :
(key == 10'b1100110101) ? 46'b0001110000101010101110100111011010000110001110 :
(key == 10'b1100110110) ? 46'b0001110000000011010100100111010111010111011101 :
(key == 10'b1100110111) ? 46'b0001101111011011111101100111010100101000111101 :
(key == 10'b1100111000) ? 46'b0001101110110100101000100111010001111010101110 :
(key == 10'b1100111001) ? 46'b0001101110001101010110100111001111001100110010 :
(key == 10'b1100111010) ? 46'b0001101101100110000111100111001100011111000111 :
(key == 10'b1100111011) ? 46'b0001101100111110111011000111001001110001110000 :
(key == 10'b1100111100) ? 46'b0001101100010111110001000111000111000100101010 :
(key == 10'b1100111101) ? 46'b0001101011110000101010000111000100010111110111 :
(key == 10'b1100111110) ? 46'b0001101011001001100110000111000001101011010101 :
(key == 10'b1100111111) ? 46'b0001101010100010100100000110111110111111000100 :
(key == 10'b1101000000) ? 46'b0001101001111011100101000110111100010011000110 :
(key == 10'b1101000001) ? 46'b0001101001010100101001000110111001100111011001 :
(key == 10'b1101000010) ? 46'b0001101000101101101111100110110110111011111101 :
(key == 10'b1101000011) ? 46'b0001101000000110111000100110110100010000110101 :
(key == 10'b1101000100) ? 46'b0001100111100000000100000110110001100101111101 :
(key == 10'b1101000101) ? 46'b0001100110111001010010100110101110111011011000 :
(key == 10'b1101000110) ? 46'b0001100110010010100011100110101100010001000100 :
(key == 10'b1101000111) ? 46'b0001100101101011110111100110101001100111000001 :
(key == 10'b1101001000) ? 46'b0001100101000101001101100110100110111101001111 :
(key == 10'b1101001001) ? 46'b0001100100011110100110100110100100010011101111 :
(key == 10'b1101001010) ? 46'b0001100011111000000010100110100001101010100001 :
(key == 10'b1101001011) ? 46'b0001100011010001100001000110011111000001100011 :
(key == 10'b1101001100) ? 46'b0001100010101011000010000110011100011000111001 :
(key == 10'b1101001101) ? 46'b0001100010000100100101100110011001110000011110 :
(key == 10'b1101001110) ? 46'b0001100001011110001011100110010111001000010101 :
(key == 10'b1101001111) ? 46'b0001100000110111110100100110010100100000011101 :
(key == 10'b1101010000) ? 46'b0001100000010001100000000110010001111000110111 :
(key == 10'b1101010001) ? 46'b0001011111101011001110000110001111010001100000 :
(key == 10'b1101010010) ? 46'b0001011111000100111111000110001100101010011101 :
(key == 10'b1101010011) ? 46'b0001011110011110110010000110001010000011101001 :
(key == 10'b1101010100) ? 46'b0001011101111000101000000110000111011101000110 :
(key == 10'b1101010101) ? 46'b0001011101010010100000100110000100110110110110 :
(key == 10'b1101010110) ? 46'b0001011100101100011011100110000010010000110110 :
(key == 10'b1101010111) ? 46'b0001011100000110011001100101111111101011000111 :
(key == 10'b1101011000) ? 46'b0001011011100000011010000101111101000101101000 :
(key == 10'b1101011001) ? 46'b0001011010111010011101000101111010100000011100 :
(key == 10'b1101011010) ? 46'b0001011010010100100010000101110111111011011110 :
(key == 10'b1101011011) ? 46'b0001011001101110101010000101110101010110110011 :
(key == 10'b1101011100) ? 46'b0001011001001000110101000101110010110010011000 :
(key == 10'b1101011101) ? 46'b0001011000100011000010000101110000001110001110 :
(key == 10'b1101011110) ? 46'b0001010111111101010010000101101101101010010100 :
(key == 10'b1101011111) ? 46'b0001010111010111100100000101101011000110101011 :
(key == 10'b1101100000) ? 46'b0001010110110001111001100101101000100011010010 :
(key == 10'b1101100001) ? 46'b0001010110001100010000100101100110000000001100 :
(key == 10'b1101100010) ? 46'b0001010101100110101010100101100011011101010011 :
(key == 10'b1101100011) ? 46'b0001010101000001000111000101100000111010101110 :
(key == 10'b1101100100) ? 46'b0001010100011011100110100101011110011000011000 :
(key == 10'b1101100101) ? 46'b0001010011110110001000000101011011110110010011 :
(key == 10'b1101100110) ? 46'b0001010011010000101100000101011001010100011100 :
(key == 10'b1101100111) ? 46'b0001010010101011010011000101010110110010111000 :
(key == 10'b1101101000) ? 46'b0001010010000101111100000101010100010001100100 :
(key == 10'b1101101001) ? 46'b0001010001100000100111100101010001110000100000 :
(key == 10'b1101101010) ? 46'b0001010000111011010110000101001111001111101100 :
(key == 10'b1101101011) ? 46'b0001010000010110000110100101001100101111001000 :
(key == 10'b1101101100) ? 46'b0001001111110000111010000101001010001110110101 :
(key == 10'b1101101101) ? 46'b0001001111001011101111100101000111101110110010 :
(key == 10'b1101101110) ? 46'b0001001110100110101000000101000101001110111110 :
(key == 10'b1101101111) ? 46'b0001001110000001100010100101000010101111011100 :
(key == 10'b1101110000) ? 46'b0001001101011100100000000101000000010000001001 :
(key == 10'b1101110001) ? 46'b0001001100110111100000000100111101110001000110 :
(key == 10'b1101110010) ? 46'b0001001100010010100010000100111011010010010011 :
(key == 10'b1101110011) ? 46'b0001001011101101100110100100111000110011110001 :
(key == 10'b1101110100) ? 46'b0001001011001000101110000100110110010101011110 :
(key == 10'b1101110101) ? 46'b0001001010100011110111100100110011110111011100 :
(key == 10'b1101110110) ? 46'b0001001001111111000011100100110001011001101001 :
(key == 10'b1101110111) ? 46'b0001001001011010010010100100101110111100000101 :
(key == 10'b1101111000) ? 46'b0001001000110101100011100100101100011110110010 :
(key == 10'b1101111001) ? 46'b0001001000010000110111000100101010000001101110 :
(key == 10'b1101111010) ? 46'b0001000111101100001101000100100111100100111011 :
(key == 10'b1101111011) ? 46'b0001000111000111100101000100100101001000010110 :
(key == 10'b1101111100) ? 46'b0001000110100011000000000100100010101100000001 :
(key == 10'b1101111101) ? 46'b0001000101111110011101100100100000001111111100 :
(key == 10'b1101111110) ? 46'b0001000101011001111101100100011101110100000111 :
(key == 10'b1101111111) ? 46'b0001000100110101011111100100011011011000100010 :
(key == 10'b1110000000) ? 46'b0001000100010001000100000100011000111101001101 :
(key == 10'b1110000001) ? 46'b0001000011101100101011000100010110100010000101 :
(key == 10'b1110000010) ? 46'b0001000011001000010100100100010100000111001101 :
(key == 10'b1110000011) ? 46'b0001000010100100000000100100010001101100101000 :
(key == 10'b1110000100) ? 46'b0001000001111111101110100100001111010010001111 :
(key == 10'b1110000101) ? 46'b0001000001011011011111100100001100111000000101 :
(key == 10'b1110000110) ? 46'b0001000000110111010010100100001010011110001100 :
(key == 10'b1110000111) ? 46'b0001000000010011001000000100001000000100100011 :
(key == 10'b1110001000) ? 46'b0000111111101111000000000100000101101011001000 :
(key == 10'b1110001001) ? 46'b0000111111001010111010000100000011010001111100 :
(key == 10'b1110001010) ? 46'b0000111110100110110111000100000000111001000000 :
(key == 10'b1110001011) ? 46'b0000111110000010110110000011111110100000010010 :
(key == 10'b1110001100) ? 46'b0000111101011110110111100011111100000111110101 :
(key == 10'b1110001101) ? 46'b0000111100111010111011100011111001101111100110 :
(key == 10'b1110001110) ? 46'b0000111100010111000010000011110111010111100111 :
(key == 10'b1110001111) ? 46'b0000111011110011001010100011110100111111110101 :
(key == 10'b1110010000) ? 46'b0000111011001111010101100011110010101000010100 :
(key == 10'b1110010001) ? 46'b0000111010101011100010100011110000010001000010 :
(key == 10'b1110010010) ? 46'b0000111010000111110010100011101101111001111110 :
(key == 10'b1110010011) ? 46'b0000111001100100000100100011101011100011001000 :
(key == 10'b1110010100) ? 46'b0000111001000000011001000011101001001100100010 :
(key == 10'b1110010101) ? 46'b0000111000011100101111100011100110110110001011 :
(key == 10'b1110010110) ? 46'b0000110111111001001001000011100100100000000100 :
(key == 10'b1110010111) ? 46'b0000110111010101100100100011100010001010001010 :
(key == 10'b1110011000) ? 46'b0000110110110010000010100011011111110100100000 :
(key == 10'b1110011001) ? 46'b0000110110001110100010100011011101011111000101 :
(key == 10'b1110011010) ? 46'b0000110101101011000101000011011011001001111001 :
(key == 10'b1110011011) ? 46'b0000110101000111101010000011011000110100111011 :
(key == 10'b1110011100) ? 46'b0000110100100100010001000011010110100000001010 :
(key == 10'b1110011101) ? 46'b0000110100000000111010100011010100001011101011 :
(key == 10'b1110011110) ? 46'b0000110011011101100110100011010001110111010111 :
(key == 10'b1110011111) ? 46'b0000110010111010010100100011001111100011010100 :
(key == 10'b1110100000) ? 46'b0000110010010111000101000011001101001111011111 :
(key == 10'b1110100001) ? 46'b0000110001110011110111100011001010111011111000 :
(key == 10'b1110100010) ? 46'b0000110001010000101101000011001000101000100001 :
(key == 10'b1110100011) ? 46'b0000110000101101100100000011000110010101011000 :
(key == 10'b1110100100) ? 46'b0000110000001010011110000011000100000010011011 :
(key == 10'b1110100101) ? 46'b0000101111100111011010000011000001101111101110 :
(key == 10'b1110100110) ? 46'b0000101111000100011000000010111111011101010000 :
(key == 10'b1110100111) ? 46'b0000101110100001011000100010111101001011000010 :
(key == 10'b1110101000) ? 46'b0000101101111110011011100010111010111000111110 :
(key == 10'b1110101001) ? 46'b0000101101011011100000100010111000100111001011 :
(key == 10'b1110101010) ? 46'b0000101100111000101000000010110110010101100110 :
(key == 10'b1110101011) ? 46'b0000101100010101110001100010110100000100010000 :
(key == 10'b1110101100) ? 46'b0000101011110010111101100010110001110011000111 :
(key == 10'b1110101101) ? 46'b0000101011010000001100000010101111100010001011 :
(key == 10'b1110101110) ? 46'b0000101010101101011100000010101101010001100001 :
(key == 10'b1110101111) ? 46'b0000101010001010101111000010101011000001000001 :
(key == 10'b1110110000) ? 46'b0000101001101000000100000010101000110000110010 :
(key == 10'b1110110001) ? 46'b0000101001000101011011000010100110100000101111 :
(key == 10'b1110110010) ? 46'b0000101000100010110100100010100100010000111100 :
(key == 10'b1110110011) ? 46'b0000101000000000010000100010100010000001010100 :
(key == 10'b1110110100) ? 46'b0000100111011101101110100010011111110001111100 :
(key == 10'b1110110101) ? 46'b0000100110111011001110100010011101100010110010 :
(key == 10'b1110110110) ? 46'b0000100110011000110001000010011011010011110110 :
(key == 10'b1110110111) ? 46'b0000100101110110010101100010011001000101001000 :
(key == 10'b1110111000) ? 46'b0000100101010011111100100010010110110110101000 :
(key == 10'b1110111001) ? 46'b0000100100110001100110000010010100101000010100 :
(key == 10'b1110111010) ? 46'b0000100100001111010001000010010010011010001111 :
(key == 10'b1110111011) ? 46'b0000100011101100111110100010010000001100011001 :
(key == 10'b1110111100) ? 46'b0000100011001010101110100010001101111110110000 :
(key == 10'b1110111101) ? 46'b0000100010101000100000100010001011110001010100 :
(key == 10'b1110111110) ? 46'b0000100010000110010100100010001001100100000111 :
(key == 10'b1110111111) ? 46'b0000100001100100001011000010000111010111000110 :
(key == 10'b1111000000) ? 46'b0000100001000010000100000010000101001010010011 :
(key == 10'b1111000001) ? 46'b0000100000011111111110100010000010111101101110 :
(key == 10'b1111000010) ? 46'b0000011111111101111011100010000000110001010110 :
(key == 10'b1111000011) ? 46'b0000011111011011111011000001111110100101001101 :
(key == 10'b1111000100) ? 46'b0000011110111001111100100001111100011001010001 :
(key == 10'b1111000101) ? 46'b0000011110011000000000000001111010001101100001 :
(key == 10'b1111000110) ? 46'b0000011101110110000101100001111000000010000000 :
(key == 10'b1111000111) ? 46'b0000011101010100001101100001110101110110101100 :
(key == 10'b1111001000) ? 46'b0000011100110010011000000001110011101011100111 :
(key == 10'b1111001001) ? 46'b0000011100010000100100100001110001100000101100 :
(key == 10'b1111001010) ? 46'b0000011011101110110010100001101111010110000010 :
(key == 10'b1111001011) ? 46'b0000011011001101000011100001101101001011100010 :
(key == 10'b1111001100) ? 46'b0000011010101011010110000001101011000001010010 :
(key == 10'b1111001101) ? 46'b0000011010001001101011000001101000110111001110 :
(key == 10'b1111001110) ? 46'b0000011001101000000010000001100110101101010110 :
(key == 10'b1111001111) ? 46'b0000011001000110011011100001100100100011101110 :
(key == 10'b1111010000) ? 46'b0000011000100100110111000001100010011010010001 :
(key == 10'b1111010001) ? 46'b0000011000000011010100100001100000010001000100 :
(key == 10'b1111010010) ? 46'b0000010111100001110100100001011110001000000001 :
(key == 10'b1111010011) ? 46'b0000010111000000010110000001011011111111001100 :
(key == 10'b1111010100) ? 46'b0000010110011110111010000001011001110110100101 :
(key == 10'b1111010101) ? 46'b0000010101111101100000100001010111101110001011 :
(key == 10'b1111010110) ? 46'b0000010101011100001000100001010101100101111100 :
(key == 10'b1111010111) ? 46'b0000010100111010110011000001010011011101111100 :
(key == 10'b1111011000) ? 46'b0000010100011001011111100001010001010110001000 :
(key == 10'b1111011001) ? 46'b0000010011111000001110000001001111001110100011 :
(key == 10'b1111011010) ? 46'b0000010011010110111111000001001101000111001000 :
(key == 10'b1111011011) ? 46'b0000010010110101110010000001001010111111111100 :
(key == 10'b1111011100) ? 46'b0000010010010100100111000001001000111000111100 :
(key == 10'b1111011101) ? 46'b0000010001110011011110000001000110110010001011 :
(key == 10'b1111011110) ? 46'b0000010001010010010111100001000100101011100100 :
(key == 10'b1111011111) ? 46'b0000010000110001010010100001000010100101001011 :
(key == 10'b1111100000) ? 46'b0000010000010000010000000001000000011110111111 :
(key == 10'b1111100001) ? 46'b0000001111101111001111100000111110011000111111 :
(key == 10'b1111100010) ? 46'b0000001111001110010001000000111100010011001100 :
(key == 10'b1111100011) ? 46'b0000001110101101010101000000111010001101100111 :
(key == 10'b1111100100) ? 46'b0000001110001100011010100000111000001000001110 :
(key == 10'b1111100101) ? 46'b0000001101101011100010100000110110000011000000 :
(key == 10'b1111100110) ? 46'b0000001101001010101100100000110011111110000000 :
(key == 10'b1111100111) ? 46'b0000001100101001111000100000110001111001001110 :
(key == 10'b1111101000) ? 46'b0000001100001001000110100000101111110100100110 :
(key == 10'b1111101001) ? 46'b0000001011101000010110100000101101110000001011 :
(key == 10'b1111101010) ? 46'b0000001011000111101001000000101011101011111110 :
(key == 10'b1111101011) ? 46'b0000001010100110111101000000101001100111111110 :
(key == 10'b1111101100) ? 46'b0000001010000110010011100000100111100100000111 :
(key == 10'b1111101101) ? 46'b0000001001100101101100000000100101100000011111 :
(key == 10'b1111101110) ? 46'b0000001001000101000110100000100011011101000011 :
(key == 10'b1111101111) ? 46'b0000001000100100100011000000100001011001110011 :
(key == 10'b1111110000) ? 46'b0000001000000100000010000000011111010110110010 :
(key == 10'b1111110001) ? 46'b0000000111100011100010100000011101010011111011 :
(key == 10'b1111110010) ? 46'b0000000111000011000101000000011011010001001111 :
(key == 10'b1111110011) ? 46'b0000000110100010101010000000011001001110110010 :
(key == 10'b1111110100) ? 46'b0000000110000010010000100000010111001100100010 :
(key == 10'b1111110101) ? 46'b0000000101100001111001100000010101001010011011 :
(key == 10'b1111110110) ? 46'b0000000101000001100100100000010011001000100010 :
(key == 10'b1111110111) ? 46'b0000000100100001010001000000010001000110110110 :
(key == 10'b1111111000) ? 46'b0000000100000001000000000000001111000101010011 :
(key == 10'b1111111001) ? 46'b0000000011100000110001000000001101000011111111 :
(key == 10'b1111111010) ? 46'b0000000011000000100100000000001011000010110111 :
(key == 10'b1111111011) ? 46'b0000000010100000011001000000001001000001111011 :
(key == 10'b1111111100) ? 46'b0000000010000000010000000000000111000001001011 :
(key == 10'b1111111101) ? 46'b0000000001100000001001000000000101000000100111 :
(key == 10'b1111111110) ? 46'b0000000001000000000100000000000011000000001111 :
(key == 10'b1111111111) ? 46'b0000000000100000000001000000000001000000000011 : 46'd0;

endmodule

`default_nettype wire
