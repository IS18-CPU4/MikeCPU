`default_nettype none

module finv
   ( input wire [31:0] x,
     output wire [31:0] y,
     output wire ovf);

   /* TODO: assumptions
    * - inputs and output are not unnormal numbers or NaN or +-inf 
    * - if e is 0, the number is interpreted as +0
    * - overflow and underflow are treated as the same for ovf wire
    * - when underflow, y will be 0
    */

   // split sequence to each subsequence
   wire xs;
   wire [7:0] xe;
   wire [22:0] xm;
   assign {xs, xe, xm} = x;

   // calc s
   wire s;
   assign s = xs;

   // calc e
   wire [7:0] e;
   assign e = (xm == 23'd0) ? 8'd254 - xe : 8'd253 - xe; 

   // calc m
   wire [22:0] m;
   wire [45:0] val;
   wire [9:0] key;
   wire [12:0] var;
   assign {key, var} = xm;
   lookup_table(key, val);
   wire [23:0] constant;
   wire [22:0] grad;
   assign {constant, grad} = {1'b1, val};
   wire [37:0] tmp_grad;
   assign tmp_grad = var * grad;
   wire [23:0] tmp_tmp_grad;
   assign tmp_tmp_grad = {10'd0, tmp_grad[37:24]};
   wire [23:0] tmp_m;
   assign tmp_m = constant - tmp_tmp_grad;
   assign m = (xm == 23'd0) ? 23'd0 : tmp_m[22:0];

   assign y = {s, e, m};

endmodule

module lookup_table
   ( input wire [9:0] key,
     output wire [45:0] value);

   assign value =
(key == 10'b0000000000) ? 46'b1111111101000000000000001111111110000000001010 :
(key == 10'b0000000001) ? 46'b1111111001000000000000001111111010000000111010 :
(key == 10'b0000000010) ? 46'b1111110101000000000000001111110110000010011001 :
(key == 10'b0000000011) ? 46'b1111110001000000000000001111110010000100101000 :
(key == 10'b0000000100) ? 46'b1111101101000000000000001111101110000111100111 :
(key == 10'b0000000101) ? 46'b1111101001010000000000001111101010001011010100 :
(key == 10'b0000000110) ? 46'b1111100101010000000000001111100110001111110001 :
(key == 10'b0000000111) ? 46'b1111100001100000000000001111100010010100111100 :
(key == 10'b0000001000) ? 46'b1111011101100000000000001111011110011010110110 :
(key == 10'b0000001001) ? 46'b1111011001010000000000001111011010100001011111 :
(key == 10'b0000001010) ? 46'b1111010101110000000000001111010110101000110110 :
(key == 10'b0000001011) ? 46'b1111010001110000000000001111010010110000111010 :
(key == 10'b0000001100) ? 46'b1111001101110000000000001111001110111001101110 :
(key == 10'b0000001101) ? 46'b1111001010000000000000001111001011000011001110 :
(key == 10'b0000001110) ? 46'b1111000110010000000000001111000111001101011100 :
(key == 10'b0000001111) ? 46'b1111000010010000000000001111000011011000011000 :
(key == 10'b0000010000) ? 46'b1110111110100000000000001110111111100100000000 :
(key == 10'b0000010001) ? 46'b1110111011000000000000001110111011110000010101 :
(key == 10'b0000010010) ? 46'b1110110110110000000000001110110111111101011000 :
(key == 10'b0000010011) ? 46'b1110110011010000000000001110110100001011000111 :
(key == 10'b0000010100) ? 46'b1110101111010000000000001110110000011001100011 :
(key == 10'b0000010101) ? 46'b1110101011100000000000001110101100101000101011 :
(key == 10'b0000010110) ? 46'b1110101000000000000000001110101000111000011111 :
(key == 10'b0000010111) ? 46'b1110100100000000000000001110100101001001000000 :
(key == 10'b0000011000) ? 46'b1110100000100000000000001110100001011010001011 :
(key == 10'b0000011001) ? 46'b1110011100110000000000001110011101101100000011 :
(key == 10'b0000011010) ? 46'b1110011001010000000000001110011001111110100110 :
(key == 10'b0000011011) ? 46'b1110010101010000000000001110010110010001110100 :
(key == 10'b0000011100) ? 46'b1110010001100000000000001110010010100101101110 :
(key == 10'b0000011101) ? 46'b1110001110000000000000001110001110111010010011 :
(key == 10'b0000011110) ? 46'b1110001010010000000000001110001011001111100010 :
(key == 10'b0000011111) ? 46'b1110000110110000000000001110000111100101011101 :
(key == 10'b0000100000) ? 46'b1110000011000000000000001110000011111100000010 :
(key == 10'b0000100001) ? 46'b1101111111100000000000001110000000010011010001 :
(key == 10'b0000100010) ? 46'b1101111011110000000000001101111100101011001010 :
(key == 10'b0000100011) ? 46'b1101111000010000000000001101111001000011101101 :
(key == 10'b0000100100) ? 46'b1101110100100000000000001101110101011100111011 :
(key == 10'b0000100101) ? 46'b1101110001000000000000001101110001110110110010 :
(key == 10'b0000100110) ? 46'b1101101101100000000000001101101110010001010010 :
(key == 10'b0000100111) ? 46'b1101101001110000000000001101101010101100011100 :
(key == 10'b0000101000) ? 46'b1101100110010000000000001101100111001000001111 :
(key == 10'b0000101001) ? 46'b1101100010110000000000001101100011100100101011 :
(key == 10'b0000101010) ? 46'b1101011111010000000000001101100000000001110001 :
(key == 10'b0000101011) ? 46'b1101011011100000000000001101011100011111011111 :
(key == 10'b0000101100) ? 46'b1101011000000000000000001101011000111101110110 :
(key == 10'b0000101101) ? 46'b1101010100100000000000001101010101011100110100 :
(key == 10'b0000101110) ? 46'b1101010001000000000000001101010001111100011100 :
(key == 10'b0000101111) ? 46'b1101001101100000000000001101001110011100101100 :
(key == 10'b0000110000) ? 46'b1101001010000000000000001101001010111101100100 :
(key == 10'b0000110001) ? 46'b1101000110100000000000001101000111011111000100 :
(key == 10'b0000110010) ? 46'b1101000011000000000000001101000100000001001011 :
(key == 10'b0000110011) ? 46'b1101000000000000000000001101000000100011111001 :
(key == 10'b0000110100) ? 46'b1100111100010000000000001100111101000111010000 :
(key == 10'b0000110101) ? 46'b1100111000110000000000001100111001101011001110 :
(key == 10'b0000110110) ? 46'b1100110101010000000000001100110110001111110011 :
(key == 10'b0000110111) ? 46'b1100110010000000000000001100110010110100111111 :
(key == 10'b0000111000) ? 46'b1100101110100000000000001100101111011010110010 :
(key == 10'b0000111001) ? 46'b1100101011010000000000001100101100000001001011 :
(key == 10'b0000111010) ? 46'b1100100111110000000000001100101000101000001010 :
(key == 10'b0000111011) ? 46'b1100100100010000000000001100100101001111110001 :
(key == 10'b0000111100) ? 46'b1100100001010000000000001100100001110111111110 :
(key == 10'b0000111101) ? 46'b1100011101100000000000001100011110100000110001 :
(key == 10'b0000111110) ? 46'b1100011010010000000000001100011011001010001010 :
(key == 10'b0000111111) ? 46'b1100010111000000000000001100010111110100001000 :
(key == 10'b0001000000) ? 46'b1100010011110000000000001100010100011110101101 :
(key == 10'b0001000001) ? 46'b1100010000010000000000001100010001001001110111 :
(key == 10'b0001000010) ? 46'b1100001100110000000000001100001101110101100111 :
(key == 10'b0001000011) ? 46'b1100001001110000000000001100001010100001111100 :
(key == 10'b0001000100) ? 46'b1100000110100000000000001100000111001110110110 :
(key == 10'b0001000101) ? 46'b1100000011010000000000001100000011111100010101 :
(key == 10'b0001000110) ? 46'b1100000000000000000000001100000000101010011001 :
(key == 10'b0001000111) ? 46'b1011111100100000000000001011111101011001000010 :
(key == 10'b0001001000) ? 46'b1011111001000000000000001011111010001000010000 :
(key == 10'b0001001001) ? 46'b1011110101110000000000001011110110111000000010 :
(key == 10'b0001001010) ? 46'b1011110010100000000000001011110011101000011000 :
(key == 10'b0001001011) ? 46'b1011101111110000000000001011110000011001010010 :
(key == 10'b0001001100) ? 46'b1011101100010000000000001011101101001010110001 :
(key == 10'b0001001101) ? 46'b1011101001000000000000001011101001111100110100 :
(key == 10'b0001001110) ? 46'b1011100110000000000000001011100110101111011010 :
(key == 10'b0001001111) ? 46'b1011100010110000000000001011100011100010100101 :
(key == 10'b0001010000) ? 46'b1011011111110000000000001011100000010110010010 :
(key == 10'b0001010001) ? 46'b1011011100100000000000001011011101001010100011 :
(key == 10'b0001010010) ? 46'b1011011001000000000000001011011001111111011001 :
(key == 10'b0001010011) ? 46'b1011010110000000000000001011010110110100110000 :
(key == 10'b0001010100) ? 46'b1011010011000000000000001011010011101010101011 :
(key == 10'b0001010101) ? 46'b1011001111110000000000001011010000100001001001 :
(key == 10'b0001010110) ? 46'b1011001100110000000000001011001101011000001010 :
(key == 10'b0001010111) ? 46'b1011001001010000000000001011001010001111101110 :
(key == 10'b0001011000) ? 46'b1011000110010000000000001011000111000111110011 :
(key == 10'b0001011001) ? 46'b1011000011010000000000001011000100000000011100 :
(key == 10'b0001011010) ? 46'b1011000000000000000000001011000000111001100110 :
(key == 10'b0001011011) ? 46'b1010111101000000000000001010111101110011010011 :
(key == 10'b0001011100) ? 46'b1010111010000000000000001010111010101101100010 :
(key == 10'b0001011101) ? 46'b1010110110110000000000001010110111101000010100 :
(key == 10'b0001011110) ? 46'b1010110100000000000000001010110100100011100110 :
(key == 10'b0001011111) ? 46'b1010110000110000000000001010110001011111011011 :
(key == 10'b0001100000) ? 46'b1010101101110000000000001010101110011011110001 :
(key == 10'b0001100001) ? 46'b1010101010100000000000001010101011011000101001 :
(key == 10'b0001100010) ? 46'b1010100111110000000000001010101000010110000010 :
(key == 10'b0001100011) ? 46'b1010100100110000000000001010100101010011111100 :
(key == 10'b0001100100) ? 46'b1010100001110000000000001010100010010010011000 :
(key == 10'b0001100101) ? 46'b1010011110100000000000001010011111010001010100 :
(key == 10'b0001100110) ? 46'b1010011011100000000000001010011100010000110010 :
(key == 10'b0001100111) ? 46'b1010011000010000000000001010011001010000110000 :
(key == 10'b0001101000) ? 46'b1010010101110000000000001010010110010001001110 :
(key == 10'b0001101001) ? 46'b1010010010110000000000001010010011010010001110 :
(key == 10'b0001101010) ? 46'b1010001111100000000000001010010000010011101110 :
(key == 10'b0001101011) ? 46'b1010001100110000000000001010001101010101101101 :
(key == 10'b0001101100) ? 46'b1010001001110000000000001010001010011000001101 :
(key == 10'b0001101101) ? 46'b1010000110110000000000001010000111011011001110 :
(key == 10'b0001101110) ? 46'b1010000011100000000000001010000100011110101111 :
(key == 10'b0001101111) ? 46'b1010000001000000000000001010000001100010101110 :
(key == 10'b0001110000) ? 46'b1001111110000000000000001001111110100111001110 :
(key == 10'b0001110001) ? 46'b1001111011000000000000001001111011101100001110 :
(key == 10'b0001110010) ? 46'b1001111000000000000000001001111000110001101101 :
(key == 10'b0001110011) ? 46'b1001110101010000000000001001110101110111101011 :
(key == 10'b0001110100) ? 46'b1001110010010000000000001001110010111110001001 :
(key == 10'b0001110101) ? 46'b1001101111010000000000001001110000000101000110 :
(key == 10'b0001110110) ? 46'b1001101100100000000000001001101101001100100011 :
(key == 10'b0001110111) ? 46'b1001101001110000000000001001101010010100011101 :
(key == 10'b0001111000) ? 46'b1001100111000000000000001001100111011100110111 :
(key == 10'b0001111001) ? 46'b1001100100000000000000001001100100100101101111 :
(key == 10'b0001111010) ? 46'b1001100001000000000000001001100001101111000111 :
(key == 10'b0001111011) ? 46'b1001011110010000000000001001011110111000111100 :
(key == 10'b0001111100) ? 46'b1001011011010000000000001001011100000011010001 :
(key == 10'b0001111101) ? 46'b1001011000100000000000001001011001001110000100 :
(key == 10'b0001111110) ? 46'b1001010101110000000000001001010110011001010100 :
(key == 10'b0001111111) ? 46'b1001010011000000000000001001010011100101000011 :
(key == 10'b0010000000) ? 46'b1001010000000000000000001001010000110001010001 :
(key == 10'b0010000001) ? 46'b1001001101010000000000001001001101111101111011 :
(key == 10'b0010000010) ? 46'b1001001010100000000000001001001011001011000100 :
(key == 10'b0010000011) ? 46'b1001000111110000000000001001001000011000101010 :
(key == 10'b0010000100) ? 46'b1001000100110000000000001001000101100110101110 :
(key == 10'b0010000101) ? 46'b1001000010010000000000001001000010110101010000 :
(key == 10'b0010000110) ? 46'b1000111111100000000000001001000000000100001111 :
(key == 10'b0010000111) ? 46'b1000111100110000000000001000111101010011101011 :
(key == 10'b0010001000) ? 46'b1000111001110000000000001000111010100011100101 :
(key == 10'b0010001001) ? 46'b1000110111010000000000001000110111110011111011 :
(key == 10'b0010001010) ? 46'b1000110100100000000000001000110101000100101111 :
(key == 10'b0010001011) ? 46'b1000110001110000000000001000110010010101111111 :
(key == 10'b0010001100) ? 46'b1000101111000000000000001000101111100111101100 :
(key == 10'b0010001101) ? 46'b1000101100010000000000001000101100111001110110 :
(key == 10'b0010001110) ? 46'b1000101001100000000000001000101010001100011101 :
(key == 10'b0010001111) ? 46'b1000100110110000000000001000100111011111100000 :
(key == 10'b0010010000) ? 46'b1000100100010000000000001000100100110010111111 :
(key == 10'b0010010001) ? 46'b1000100001100000000000001000100010000110111011 :
(key == 10'b0010010010) ? 46'b1000011110110000000000001000011111011011010011 :
(key == 10'b0010010011) ? 46'b1000011100010000000000001000011100110000000110 :
(key == 10'b0010010100) ? 46'b1000011001100000000000001000011010000101010111 :
(key == 10'b0010010101) ? 46'b1000010110110000000000001000010111011011000011 :
(key == 10'b0010010110) ? 46'b1000010100010000000000001000010100110001001010 :
(key == 10'b0010010111) ? 46'b1000010001100000000000001000010010000111101110 :
(key == 10'b0010011000) ? 46'b1000001111000000000000001000001111011110101101 :
(key == 10'b0010011001) ? 46'b1000001100010000000000001000001100110110001000 :
(key == 10'b0010011010) ? 46'b1000001001100000000000001000001010001101111111 :
(key == 10'b0010011011) ? 46'b1000000110110000000000001000000111100110010000 :
(key == 10'b0010011100) ? 46'b1000000100010000000000001000000100111110111101 :
(key == 10'b0010011101) ? 46'b1000000001110000000000001000000010011000000101 :
(key == 10'b0010011110) ? 46'b0111111111010000000000000111111111110001101000 :
(key == 10'b0010011111) ? 46'b0111111100100000000000000111111101001011100110 :
(key == 10'b0010100000) ? 46'b0111111010000000000000000111111010100101111111 :
(key == 10'b0010100001) ? 46'b0111110111010000000000000111111000000000110011 :
(key == 10'b0010100010) ? 46'b0111110100110000000000000111110101011100000001 :
(key == 10'b0010100011) ? 46'b0111110010010000000000000111110010110111101011 :
(key == 10'b0010100100) ? 46'b0111101111110000000000000111110000010011101110 :
(key == 10'b0010100101) ? 46'b0111101101000000000000000111101101110000001101 :
(key == 10'b0010100110) ? 46'b0111101010100000000000000111101011001101000101 :
(key == 10'b0010100111) ? 46'b0111101000000000000000000111101000101010011000 :
(key == 10'b0010101000) ? 46'b0111100101100000000000000111100110001000000100 :
(key == 10'b0010101001) ? 46'b0111100010110000000000000111100011100110001100 :
(key == 10'b0010101010) ? 46'b0111100000100000000000000111100001000100101101 :
(key == 10'b0010101011) ? 46'b0111011110000000000000000111011110100011101000 :
(key == 10'b0010101100) ? 46'b0111011011100000000000000111011100000010111101 :
(key == 10'b0010101101) ? 46'b0111011001000000000000000111011001100010101100 :
(key == 10'b0010101110) ? 46'b0111010110100000000000000111010111000010110011 :
(key == 10'b0010101111) ? 46'b0111010011110000000000000111010100100011010101 :
(key == 10'b0010110000) ? 46'b0111010001100000000000000111010010000100010000 :
(key == 10'b0010110001) ? 46'b0111001111000000000000000111001111100101100110 :
(key == 10'b0010110010) ? 46'b0111001100100000000000000111001101000111010011 :
(key == 10'b0010110011) ? 46'b0111001010000000000000000111001010101001011011 :
(key == 10'b0010110100) ? 46'b0111000111100000000000000111001000001011111100 :
(key == 10'b0010110101) ? 46'b0111000101010000000000000111000101101110110101 :
(key == 10'b0010110110) ? 46'b0111000010110000000000000111000011010010000111 :
(key == 10'b0010110111) ? 46'b0111000000100000000000000111000000110101110010 :
(key == 10'b0010111000) ? 46'b0110111110000000000000000110111110011001110111 :
(key == 10'b0010111001) ? 46'b0110111011100000000000000110111011111110010100 :
(key == 10'b0010111010) ? 46'b0110111001000000000000000110111001100011001010 :
(key == 10'b0010111011) ? 46'b0110110110100000000000000110110111001000011000 :
(key == 10'b0010111100) ? 46'b0110110100000000000000000110110100101101111111 :
(key == 10'b0010111101) ? 46'b0110110001100000000000000110110010010011111110 :
(key == 10'b0010111110) ? 46'b0110101111010000000000000110101111111010010110 :
(key == 10'b0010111111) ? 46'b0110101100110000000000000110101101100001000101 :
(key == 10'b0011000000) ? 46'b0110101010100000000000000110101011001000001101 :
(key == 10'b0011000001) ? 46'b0110101000000000000000000110101000101111101101 :
(key == 10'b0011000010) ? 46'b0110100101110000000000000110100110010111100101 :
(key == 10'b0011000011) ? 46'b0110100011100000000000000110100011111111110101 :
(key == 10'b0011000100) ? 46'b0110100001010000000000000110100001101000011100 :
(key == 10'b0011000101) ? 46'b0110011110100000000000000110011111010001011101 :
(key == 10'b0011000110) ? 46'b0110011100010000000000000110011100111010110100 :
(key == 10'b0011000111) ? 46'b0110011010000000000000000110011010100100100011 :
(key == 10'b0011001000) ? 46'b0110010111110000000000000110011000001110101001 :
(key == 10'b0011001001) ? 46'b0110010101100000000000000110010101111001000111 :
(key == 10'b0011001010) ? 46'b0110010010110000000000000110010011100011111101 :
(key == 10'b0011001011) ? 46'b0110010000110000000000000110010001001111001001 :
(key == 10'b0011001100) ? 46'b0110001110010000000000000110001110111010101110 :
(key == 10'b0011001101) ? 46'b0110001100000000000000000110001100100110101001 :
(key == 10'b0011001110) ? 46'b0110001001110000000000000110001010010010111011 :
(key == 10'b0011001111) ? 46'b0110000111100000000000000110000111111111100100 :
(key == 10'b0011010000) ? 46'b0110000101010000000000000110000101101100100100 :
(key == 10'b0011010001) ? 46'b0110000010110000000000000110000011011001111011 :
(key == 10'b0011010010) ? 46'b0110000000100000000000000110000001000111101001 :
(key == 10'b0011010011) ? 46'b0101111110010000000000000101111110110101101110 :
(key == 10'b0011010100) ? 46'b0101111100000000000000000101111100100100001001 :
(key == 10'b0011010101) ? 46'b0101111001110000000000000101111010010010111011 :
(key == 10'b0011010110) ? 46'b0101110111010000000000000101111000000010000100 :
(key == 10'b0011010111) ? 46'b0101110101010000000000000101110101110001100010 :
(key == 10'b0011011000) ? 46'b0101110011000000000000000101110011100001010111 :
(key == 10'b0011011001) ? 46'b0101110000110000000000000101110001010001100010 :
(key == 10'b0011011010) ? 46'b0101101110010000000000000101101111000010000100 :
(key == 10'b0011011011) ? 46'b0101101100100000000000000101101100110010111011 :
(key == 10'b0011011100) ? 46'b0101101010000000000000000101101010100100001010 :
(key == 10'b0011011101) ? 46'b0101101000000000000000000101101000010101101101 :
(key == 10'b0011011110) ? 46'b0101100101010000000000000101100110000111101000 :
(key == 10'b0011011111) ? 46'b0101100011100000000000000101100011111001110110 :
(key == 10'b0011100000) ? 46'b0101100001000000000000000101100001101100011100 :
(key == 10'b0011100001) ? 46'b0101011111000000000000000101011111011111010111 :
(key == 10'b0011100010) ? 46'b0101011100110000000000000101011101010010101000 :
(key == 10'b0011100011) ? 46'b0101011010100000000000000101011011000110001111 :
(key == 10'b0011100100) ? 46'b0101011000010000000000000101011000111010001011 :
(key == 10'b0011100101) ? 46'b0101010110010000000000000101010110101110011100 :
(key == 10'b0011100110) ? 46'b0101010100000000000000000101010100100011000011 :
(key == 10'b0011100111) ? 46'b0101010001110000000000000101010010010111111110 :
(key == 10'b0011101000) ? 46'b0101001111100000000000000101010000001101010000 :
(key == 10'b0011101001) ? 46'b0101001101100000000000000101001110000010110110 :
(key == 10'b0011101010) ? 46'b0101001011010000000000000101001011111000110010 :
(key == 10'b0011101011) ? 46'b0101001001000000000000000101001001101111000011 :
(key == 10'b0011101100) ? 46'b0101000111010000000000000101000111100101101000 :
(key == 10'b0011101101) ? 46'b0101000101000000000000000101000101011100100010 :
(key == 10'b0011101110) ? 46'b0101000010110000000000000101000011010011110001 :
(key == 10'b0011101111) ? 46'b0101000000110000000000000101000001001011010101 :
(key == 10'b0011110000) ? 46'b0100111110110000000000000100111111000011001110 :
(key == 10'b0011110001) ? 46'b0100111100100000000000000100111100111011011100 :
(key == 10'b0011110010) ? 46'b0100111010000000000000000100111010110011111110 :
(key == 10'b0011110011) ? 46'b0100111000000000000000000100111000101100110101 :
(key == 10'b0011110100) ? 46'b0100110110010000000000000100110110100101111111 :
(key == 10'b0011110101) ? 46'b0100110100000000000000000100110100011111011111 :
(key == 10'b0011110110) ? 46'b0100110010000000000000000100110010011001010010 :
(key == 10'b0011110111) ? 46'b0100101111100000000000000100110000010011011011 :
(key == 10'b0011111000) ? 46'b0100101101100000000000000100101110001101110111 :
(key == 10'b0011111001) ? 46'b0100101011110000000000000100101100001000100110 :
(key == 10'b0011111010) ? 46'b0100101001110000000000000100101010000011101011 :
(key == 10'b0011111011) ? 46'b0100100111100000000000000100100111111111000011 :
(key == 10'b0011111100) ? 46'b0100100101100000000000000100100101111010110000 :
(key == 10'b0011111101) ? 46'b0100100011010000000000000100100011110110110000 :
(key == 10'b0011111110) ? 46'b0100100001010000000000000100100001110011000100 :
(key == 10'b0011111111) ? 46'b0100011111000000000000000100011111101111101011 :
(key == 10'b0100000000) ? 46'b0100011101000000000000000100011101101100100111 :
(key == 10'b0100000001) ? 46'b0100011011000000000000000100011011101001110110 :
(key == 10'b0100000010) ? 46'b0100011001000000000000000100011001100111011001 :
(key == 10'b0100000011) ? 46'b0100010111000000000000000100010111100101001111 :
(key == 10'b0100000100) ? 46'b0100010101000000000000000100010101100011011000 :
(key == 10'b0100000101) ? 46'b0100010011000000000000000100010011100001110101 :
(key == 10'b0100000110) ? 46'b0100010001000000000000000100010001100000100101 :
(key == 10'b0100000111) ? 46'b0100001111000000000000000100001111011111101001 :
(key == 10'b0100001000) ? 46'b0100001101000000000000000100001101011110111111 :
(key == 10'b0100001001) ? 46'b0100001011000000000000000100001011011110101001 :
(key == 10'b0100001010) ? 46'b0100001001000000000000000100001001011110100110 :
(key == 10'b0100001011) ? 46'b0100000111000000000000000100000111011110110110 :
(key == 10'b0100001100) ? 46'b0100000101000000000000000100000101011111011001 :
(key == 10'b0100001101) ? 46'b0100000011000000000000000100000011100000001111 :
(key == 10'b0100001110) ? 46'b0100000001000000000000000100000001100001010111 :
(key == 10'b0100001111) ? 46'b0011111111000000000000000011111111100010110011 :
(key == 10'b0100010000) ? 46'b0011111101000000000000000011111101100100100010 :
(key == 10'b0100010001) ? 46'b0011111011010000000000000011111011100110100010 :
(key == 10'b0100010010) ? 46'b0011111001010000000000000011111001101000110110 :
(key == 10'b0100010011) ? 46'b0011110111000000000000000011110111101011011100 :
(key == 10'b0100010100) ? 46'b0011110101010000000000000011110101101110010101 :
(key == 10'b0100010101) ? 46'b0011110011010000000000000011110011110001100000 :
(key == 10'b0100010110) ? 46'b0011110001010000000000000011110001110100111101 :
(key == 10'b0100010111) ? 46'b0011101111100000000000000011101111111000101101 :
(key == 10'b0100011000) ? 46'b0011101101010000000000000011101101111100110000 :
(key == 10'b0100011001) ? 46'b0011101011100000000000000011101100000001000100 :
(key == 10'b0100011010) ? 46'b0011101001110000000000000011101010000101101010 :
(key == 10'b0100011011) ? 46'b0011100111110000000000000011101000001010100010 :
(key == 10'b0100011100) ? 46'b0011100101110000000000000011100110001111101101 :
(key == 10'b0100011101) ? 46'b0011100100000000000000000011100100010101001010 :
(key == 10'b0100011110) ? 46'b0011100010000000000000000011100010011010111000 :
(key == 10'b0100011111) ? 46'b0011100000000000000000000011100000100000111001 :
(key == 10'b0100100000) ? 46'b0011011110010000000000000011011110100111001011 :
(key == 10'b0100100001) ? 46'b0011011100010000000000000011011100101101110000 :
(key == 10'b0100100010) ? 46'b0011011010010000000000000011011010110100100110 :
(key == 10'b0100100011) ? 46'b0011011000100000000000000011011000111011101101 :
(key == 10'b0100100100) ? 46'b0011010110100000000000000011010111000011000110 :
(key == 10'b0100100101) ? 46'b0011010100100000000000000011010101001010110001 :
(key == 10'b0100100110) ? 46'b0011010010110000000000000011010011010010101101 :
(key == 10'b0100100111) ? 46'b0011010001000000000000000011010001011010111010 :
(key == 10'b0100101000) ? 46'b0011001111000000000000000011001111100011011010 :
(key == 10'b0100101001) ? 46'b0011001101010000000000000011001101101100001010 :
(key == 10'b0100101010) ? 46'b0011001011100000000000000011001011110101001100 :
(key == 10'b0100101011) ? 46'b0011001001100000000000000011001001111110011111 :
(key == 10'b0100101100) ? 46'b0011000111100000000000000011001000001000000100 :
(key == 10'b0100101101) ? 46'b0011000101110000000000000011000110010001111001 :
(key == 10'b0100101110) ? 46'b0011000100000000000000000011000100011011111111 :
(key == 10'b0100101111) ? 46'b0011000010010000000000000011000010100110010111 :
(key == 10'b0100110000) ? 46'b0011000000100000000000000011000000110000111111 :
(key == 10'b0100110001) ? 46'b0010111110100000000000000010111110111011111001 :
(key == 10'b0100110010) ? 46'b0010111100110000000000000010111101000111000011 :
(key == 10'b0100110011) ? 46'b0010111011000000000000000010111011010010011110 :
(key == 10'b0100110100) ? 46'b0010111001000000000000000010111001011110001010 :
(key == 10'b0100110101) ? 46'b0010110111010000000000000010110111101010000111 :
(key == 10'b0100110110) ? 46'b0010110101100000000000000010110101110110010100 :
(key == 10'b0100110111) ? 46'b0010110011100000000000000010110100000010110010 :
(key == 10'b0100111000) ? 46'b0010110001110000000000000010110010001111100001 :
(key == 10'b0100111001) ? 46'b0010110000000000000000000010110000011100100000 :
(key == 10'b0100111010) ? 46'b0010101110010000000000000010101110101001101111 :
(key == 10'b0100111011) ? 46'b0010101100100000000000000010101100110111010000 :
(key == 10'b0100111100) ? 46'b0010101010100000000000000010101011000101000001 :
(key == 10'b0100111101) ? 46'b0010101001000000000000000010101001010011000001 :
(key == 10'b0100111110) ? 46'b0010100111000000000000000010100111100001010010 :
(key == 10'b0100111111) ? 46'b0010100101010000000000000010100101101111110100 :
(key == 10'b0101000000) ? 46'b0010100011100000000000000010100011111110100101 :
(key == 10'b0101000001) ? 46'b0010100001110000000000000010100010001101100111 :
(key == 10'b0101000010) ? 46'b0010100000000000000000000010100000011100111001 :
(key == 10'b0101000011) ? 46'b0010011110010000000000000010011110101100011011 :
(key == 10'b0101000100) ? 46'b0010011100100000000000000010011100111100001101 :
(key == 10'b0101000101) ? 46'b0010011010110000000000000010011011001100001111 :
(key == 10'b0101000110) ? 46'b0010011001010000000000000010011001011100100000 :
(key == 10'b0101000111) ? 46'b0010010111010000000000000010010111101101000010 :
(key == 10'b0101001000) ? 46'b0010010101100000000000000010010101111101110100 :
(key == 10'b0101001001) ? 46'b0010010100000000000000000010010100001110110101 :
(key == 10'b0101001010) ? 46'b0010010010000000000000000010010010100000000110 :
(key == 10'b0101001011) ? 46'b0010010000010000000000000010010000110001100110 :
(key == 10'b0101001100) ? 46'b0010001110110000000000000010001111000011010111 :
(key == 10'b0101001101) ? 46'b0010001101000000000000000010001101010101010110 :
(key == 10'b0101001110) ? 46'b0010001011010000000000000010001011100111100110 :
(key == 10'b0101001111) ? 46'b0010001001110000000000000010001001111010000101 :
(key == 10'b0101010000) ? 46'b0010000111110000000000000010001000001100110011 :
(key == 10'b0101010001) ? 46'b0010000110000000000000000010000110011111110001 :
(key == 10'b0101010010) ? 46'b0010000100100000000000000010000100110010111110 :
(key == 10'b0101010011) ? 46'b0010000010110000000000000010000011000110011010 :
(key == 10'b0101010100) ? 46'b0010000001000000000000000010000001011010000110 :
(key == 10'b0101010101) ? 46'b0001111111010000000000000001111111101110000001 :
(key == 10'b0101010110) ? 46'b0001111101100000000000000001111110000010001011 :
(key == 10'b0101010111) ? 46'b0001111100000000000000000001111100010110100100 :
(key == 10'b0101011000) ? 46'b0001111010010000000000000001111010101011001101 :
(key == 10'b0101011001) ? 46'b0001111000100000000000000001111001000000000101 :
(key == 10'b0101011010) ? 46'b0001110111000000000000000001110111010101001011 :
(key == 10'b0101011011) ? 46'b0001110101010000000000000001110101101010100000 :
(key == 10'b0101011100) ? 46'b0001110011100000000000000001110100000000000101 :
(key == 10'b0101011101) ? 46'b0001110010000000000000000001110010010101110111 :
(key == 10'b0101011110) ? 46'b0001110000010000000000000001110000101011111001 :
(key == 10'b0101011111) ? 46'b0001101110110000000000000001101111000010001010 :
(key == 10'b0101100000) ? 46'b0001101100110000000000000001101101011000101010 :
(key == 10'b0101100001) ? 46'b0001101011100000000000000001101011101111011000 :
(key == 10'b0101100010) ? 46'b0001101001110000000000000001101010000110010101 :
(key == 10'b0101100011) ? 46'b0001101000000000000000000001101000011101100000 :
(key == 10'b0101100100) ? 46'b0001100110100000000000000001100110110100111010 :
(key == 10'b0101100101) ? 46'b0001100100110000000000000001100101001100100011 :
(key == 10'b0101100110) ? 46'b0001100011010000000000000001100011100100011010 :
(key == 10'b0101100111) ? 46'b0001100001100000000000000001100001111100011111 :
(key == 10'b0101101000) ? 46'b0001100000000000000000000001100000010100110011 :
(key == 10'b0101101001) ? 46'b0001011110010000000000000001011110101101010110 :
(key == 10'b0101101010) ? 46'b0001011100110000000000000001011101000110000110 :
(key == 10'b0101101011) ? 46'b0001011011010000000000000001011011011111000101 :
(key == 10'b0101101100) ? 46'b0001011001100000000000000001011001111000010010 :
(key == 10'b0101101101) ? 46'b0001011000000000000000000001011000010001101101 :
(key == 10'b0101101110) ? 46'b0001010110010000000000000001010110101011010111 :
(key == 10'b0101101111) ? 46'b0001010100110000000000000001010101000101001110 :
(key == 10'b0101110000) ? 46'b0001010011000000000000000001010011011111010100 :
(key == 10'b0101110001) ? 46'b0001010001100000000000000001010001111001101000 :
(key == 10'b0101110010) ? 46'b0001001111110000000000000001010000010100001010 :
(key == 10'b0101110011) ? 46'b0001001110100000000000000001001110101110111001 :
(key == 10'b0101110100) ? 46'b0001001100110000000000000001001101001001110111 :
(key == 10'b0101110101) ? 46'b0001001011000000000000000001001011100101000010 :
(key == 10'b0101110110) ? 46'b0001001001100000000000000001001010000000011100 :
(key == 10'b0101110111) ? 46'b0001001000000000000000000001001000011100000011 :
(key == 10'b0101111000) ? 46'b0001000110100000000000000001000110110111111000 :
(key == 10'b0101111001) ? 46'b0001000100110000000000000001000101010011111010 :
(key == 10'b0101111010) ? 46'b0001000011010000000000000001000011110000001011 :
(key == 10'b0101111011) ? 46'b0001000001110000000000000001000010001100101000 :
(key == 10'b0101111100) ? 46'b0001000000010000000000000001000000101001010011 :
(key == 10'b0101111101) ? 46'b0000111110110000000000000000111111000110001101 :
(key == 10'b0101111110) ? 46'b0000111101010000000000000000111101100011010011 :
(key == 10'b0101111111) ? 46'b0000111011100000000000000000111100000000101000 :
(key == 10'b0110000000) ? 46'b0000111010000000000000000000111010011110001001 :
(key == 10'b0110000001) ? 46'b0000111000110000000000000000111000111011111000 :
(key == 10'b0110000010) ? 46'b0000110111000000000000000000110111011001110100 :
(key == 10'b0110000011) ? 46'b0000110101010000000000000000110101110111111110 :
(key == 10'b0110000100) ? 46'b0000110011110000000000000000110100010110010101 :
(key == 10'b0110000101) ? 46'b0000110010100000000000000000110010110100111001 :
(key == 10'b0110000110) ? 46'b0000110000110000000000000000110001010011101011 :
(key == 10'b0110000111) ? 46'b0000101111100000000000000000101111110010101001 :
(key == 10'b0110001000) ? 46'b0000101110000000000000000000101110010001110101 :
(key == 10'b0110001001) ? 46'b0000101100010000000000000000101100110001001110 :
(key == 10'b0110001010) ? 46'b0000101010110000000000000000101011010000110100 :
(key == 10'b0110001011) ? 46'b0000101001100000000000000000101001110000100110 :
(key == 10'b0110001100) ? 46'b0000101000000000000000000000101000010000100110 :
(key == 10'b0110001101) ? 46'b0000100110100000000000000000100110110000110011 :
(key == 10'b0110001110) ? 46'b0000100101000000000000000000100101010001001101 :
(key == 10'b0110001111) ? 46'b0000100011100000000000000000100011110001110100 :
(key == 10'b0110010000) ? 46'b0000100001110000000000000000100010010010101000 :
(key == 10'b0110010001) ? 46'b0000100000100000000000000000100000110011100111 :
(key == 10'b0110010010) ? 46'b0000011110110000000000000000011111010100110101 :
(key == 10'b0110010011) ? 46'b0000011101100000000000000000011101110110001111 :
(key == 10'b0110010100) ? 46'b0000011100010000000000000000011100010111110101 :
(key == 10'b0110010101) ? 46'b0000011010100000000000000000011010111001101001 :
(key == 10'b0110010110) ? 46'b0000011001000000000000000000011001011011101001 :
(key == 10'b0110010111) ? 46'b0000010111100000000000000000010111111101110101 :
(key == 10'b0110011000) ? 46'b0000010110010000000000000000010110100000001110 :
(key == 10'b0110011001) ? 46'b0000010100110000000000000000010101000010110100 :
(key == 10'b0110011010) ? 46'b0000010011000000000000000000010011100101100110 :
(key == 10'b0110011011) ? 46'b0000010001110000000000000000010010001000100101 :
(key == 10'b0110011100) ? 46'b0000010000100000000000000000010000101011101111 :
(key == 10'b0110011101) ? 46'b0000001110110000000000000000001111001111000111 :
(key == 10'b0110011110) ? 46'b0000001101010000000000000000001101110010101011 :
(key == 10'b0110011111) ? 46'b0000001100000000000000000000001100010110011011 :
(key == 10'b0110100000) ? 46'b0000001010100000000000000000001010111010010111 :
(key == 10'b0110100001) ? 46'b0000001001000000000000000000001001011110100001 :
(key == 10'b0110100010) ? 46'b0000000111110000000000000000001000000010110101 :
(key == 10'b0110100011) ? 46'b0000000110010000000000000000000110100111010110 :
(key == 10'b0110100100) ? 46'b0000000100110000000000000000000101001100000100 :
(key == 10'b0110100101) ? 46'b0000000011010000000000000000000011110000111101 :
(key == 10'b0110100110) ? 46'b0000000010000000000000000000000010010110000010 :
(key == 10'b0110100111) ? 46'b0000000000110000000000000000000000111011010100 :
(key == 10'b0110101000) ? 46'b1111111110100000000000001111111111000001100010 :
(key == 10'b0110101001) ? 46'b1111111011100000000000001111111100001100110110 :
(key == 10'b0110101010) ? 46'b1111111000100000000000001111111001011000100001 :
(key == 10'b0110101011) ? 46'b1111110110000000000000001111110110100100100011 :
(key == 10'b0110101100) ? 46'b1111110011100000000000001111110011110000111110 :
(key == 10'b0110101101) ? 46'b1111110000000000000000001111110000111101110000 :
(key == 10'b0110101110) ? 46'b1111101101100000000000001111101110001010111011 :
(key == 10'b0110101111) ? 46'b1111101011000000000000001111101011011000011011 :
(key == 10'b0110110000) ? 46'b1111100111100000000000001111101000100110010101 :
(key == 10'b0110110001) ? 46'b1111100101000000000000001111100101110100100110 :
(key == 10'b0110110010) ? 46'b1111100010000000000000001111100011000011001101 :
(key == 10'b0110110011) ? 46'b1111011111100000000000001111100000010010001100 :
(key == 10'b0110110100) ? 46'b1111011100100000000000001111011101100001100011 :
(key == 10'b0110110101) ? 46'b1111011010000000000000001111011010110001010000 :
(key == 10'b0110110110) ? 46'b1111010111100000000000001111011000000001010100 :
(key == 10'b0110110111) ? 46'b1111010100100000000000001111010101010001110001 :
(key == 10'b0110111000) ? 46'b1111010010000000000000001111010010100010100011 :
(key == 10'b0110111001) ? 46'b1111001110100000000000001111001111110011101110 :
(key == 10'b0110111010) ? 46'b1111001100100000000000001111001101000101001111 :
(key == 10'b0110111011) ? 46'b1111001001100000000000001111001010010111000110 :
(key == 10'b0110111100) ? 46'b1111000111000000000000001111000111101001010100 :
(key == 10'b0110111101) ? 46'b1111000100000000000000001111000100111011111001 :
(key == 10'b0110111110) ? 46'b1111000001100000000000001111000010001110110100 :
(key == 10'b0110111111) ? 46'b1110111111000000000000001110111111100010000111 :
(key == 10'b0111000000) ? 46'b1110111100000000000000001110111100110101101111 :
(key == 10'b0111000001) ? 46'b1110111001100000000000001110111010001001101111 :
(key == 10'b0111000010) ? 46'b1110110110100000000000001110110111011110000100 :
(key == 10'b0111000011) ? 46'b1110110100100000000000001110110100110010110000 :
(key == 10'b0111000100) ? 46'b1110110001100000000000001110110010000111110011 :
(key == 10'b0111000101) ? 46'b1110101111000000000000001110101111011101001010 :
(key == 10'b0111000110) ? 46'b1110101100000000000000001110101100110010111001 :
(key == 10'b0111000111) ? 46'b1110101001100000000000001110101010001000111110 :
(key == 10'b0111001000) ? 46'b1110100111000000000000001110100111011111011001 :
(key == 10'b0111001001) ? 46'b1110100100000000000000001110100100110110001001 :
(key == 10'b0111001010) ? 46'b1110100001100000000000001110100010001101010000 :
(key == 10'b0111001011) ? 46'b1110011111000000000000001110011111100100101011 :
(key == 10'b0111001100) ? 46'b1110011100100000000000001110011100111100011101 :
(key == 10'b0111001101) ? 46'b1110011001100000000000001110011010010100100110 :
(key == 10'b0111001110) ? 46'b1110010111000000000000001110010111101101000100 :
(key == 10'b0111001111) ? 46'b1110010100100000000000001110010101000101110110 :
(key == 10'b0111010000) ? 46'b1110010010000000000000001110010010011110111111 :
(key == 10'b0111010001) ? 46'b1110001111100000000000001110001111111000011101 :
(key == 10'b0111010010) ? 46'b1110001100100000000000001110001101010010010001 :
(key == 10'b0111010011) ? 46'b1110001010000000000000001110001010101100011010 :
(key == 10'b0111010100) ? 46'b1110000111100000000000001110001000000110111000 :
(key == 10'b0111010101) ? 46'b1110000101000000000000001110000101100001101100 :
(key == 10'b0111010110) ? 46'b1110000010100000000000001110000010111100110101 :
(key == 10'b0111010111) ? 46'b1101111111100000000000001110000000011000010100 :
(key == 10'b0111011000) ? 46'b1101111101100000000000001101111101110100000110 :
(key == 10'b0111011001) ? 46'b1101111010100000000000001101111011010000001111 :
(key == 10'b0111011010) ? 46'b1101111000000000000000001101111000101100101100 :
(key == 10'b0111011011) ? 46'b1101110101100000000000001101110110001001011101 :
(key == 10'b0111011100) ? 46'b1101110011000000000000001101110011100110100101 :
(key == 10'b0111011101) ? 46'b1101110000000000000000001101110001000100000001 :
(key == 10'b0111011110) ? 46'b1101101110000000000000001101101110100001110001 :
(key == 10'b0111011111) ? 46'b1101101011100000000000001101101011111111110110 :
(key == 10'b0111100000) ? 46'b1101101001000000000000001101101001011110010000 :
(key == 10'b0111100001) ? 46'b1101100110000000000000001101100110111101000000 :
(key == 10'b0111100010) ? 46'b1101100011100000000000001101100100011100000011 :
(key == 10'b0111100011) ? 46'b1101100001100000000000001101100001111011011010 :
(key == 10'b0111100100) ? 46'b1101011111000000000000001101011111011011000101 :
(key == 10'b0111100101) ? 46'b1101011100000000000000001101011100111011000111 :
(key == 10'b0111100110) ? 46'b1101011010000000000000001101011010011011011011 :
(key == 10'b0111100111) ? 46'b1101010111100000000000001101010111111100000100 :
(key == 10'b0111101000) ? 46'b1101010101000000000000001101010101011101000001 :
(key == 10'b0111101001) ? 46'b1101010010000000000000001101010010111110010011 :
(key == 10'b0111101010) ? 46'b1101010000000000000000001101010000011111111001 :
(key == 10'b0111101011) ? 46'b1101001101100000000000001101001110000001110010 :
(key == 10'b0111101100) ? 46'b1101001011000000000000001101001011100011111111 :
(key == 10'b0111101101) ? 46'b1101001000100000000000001101001001000110100001 :
(key == 10'b0111101110) ? 46'b1101000110000000000000001101000110101001010111 :
(key == 10'b0111101111) ? 46'b1101000011100000000000001101000100001100100000 :
(key == 10'b0111110000) ? 46'b1101000001000000000000001101000001101111111101 :
(key == 10'b0111110001) ? 46'b1100111110100000000000001100111111010011101110 :
(key == 10'b0111110010) ? 46'b1100111100000000000000001100111100110111110011 :
(key == 10'b0111110011) ? 46'b1100111001100000000000001100111010011100001011 :
(key == 10'b0111110100) ? 46'b1100110111100000000000001100111000000000110110 :
(key == 10'b0111110101) ? 46'b1100110101000000000000001100110101100101110110 :
(key == 10'b0111110110) ? 46'b1100110010100000000000001100110011001011001000 :
(key == 10'b0111110111) ? 46'b1100110000100000000000001100110000110000101110 :
(key == 10'b0111111000) ? 46'b1100101110000000000000001100101110010110101000 :
(key == 10'b0111111001) ? 46'b1100101011000000000000001100101011111100110110 :
(key == 10'b0111111010) ? 46'b1100101001000000000000001100101001100011010110 :
(key == 10'b0111111011) ? 46'b1100100110100000000000001100100111001010001001 :
(key == 10'b0111111100) ? 46'b1100100100000000000000001100100100110001010000 :
(key == 10'b0111111101) ? 46'b1100100001100000000000001100100010011000101010 :
(key == 10'b0111111110) ? 46'b1100011111100000000000001100100000000000010110 :
(key == 10'b0111111111) ? 46'b1100011101000000000000001100011101101000010111 :
(key == 10'b1000000000) ? 46'b1100011010100000000000001100011011010000101001 :
(key == 10'b1000000001) ? 46'b1100011000000000000000001100011000111001010000 :
(key == 10'b1000000010) ? 46'b1100010110000000000000001100010110100010001000 :
(key == 10'b1000000011) ? 46'b1100010011000000000000001100010100001011010101 :
(key == 10'b1000000100) ? 46'b1100010001000000000000001100010001110100110011 :
(key == 10'b1000000101) ? 46'b1100001111000000000000001100001111011110100100 :
(key == 10'b1000000110) ? 46'b1100001100100000000000001100001101001000101000 :
(key == 10'b1000000111) ? 46'b1100001010000000000000001100001010110010111110 :
(key == 10'b1000001000) ? 46'b1100001000000000000000001100001000011101100110 :
(key == 10'b1000001001) ? 46'b1100000101100000000000001100000110001000100010 :
(key == 10'b1000001010) ? 46'b1100000011100000000000001100000011110011110000 :
(key == 10'b1000001011) ? 46'b1100000001000000000000001100000001011111010010 :
(key == 10'b1000001100) ? 46'b1011111111000000000000001011111111001011000100 :
(key == 10'b1000001101) ? 46'b1011111100100000000000001011111100110111001001 :
(key == 10'b1000001110) ? 46'b1011111010000000000000001011111010100011100001 :
(key == 10'b1000001111) ? 46'b1011110111100000000000001011111000010000001100 :
(key == 10'b1000010000) ? 46'b1011110101100000000000001011110101111101000111 :
(key == 10'b1000010001) ? 46'b1011110011000000000000001011110011101010010110 :
(key == 10'b1000010010) ? 46'b1011110001000000000000001011110001010111110110 :
(key == 10'b1000010011) ? 46'b1011101110100000000000001011101111000101101000 :
(key == 10'b1000010100) ? 46'b1011101100100000000000001011101100110011101101 :
(key == 10'b1000010101) ? 46'b1011101010000000000000001011101010100010000100 :
(key == 10'b1000010110) ? 46'b1011101000000000000000001011101000010000101100 :
(key == 10'b1000010111) ? 46'b1011100101100000000000001011100101111111100111 :
(key == 10'b1000011000) ? 46'b1011100011000000000000001011100011101110110011 :
(key == 10'b1000011001) ? 46'b1011100001000000000000001011100001011110010001 :
(key == 10'b1000011010) ? 46'b1011011111000000000000001011011111001110000000 :
(key == 10'b1000011011) ? 46'b1011011100100000000000001011011100111110000010 :
(key == 10'b1000011100) ? 46'b1011011010000000000000001011011010101110010110 :
(key == 10'b1000011101) ? 46'b1011011000000000000000001011011000011110111010 :
(key == 10'b1000011110) ? 46'b1011010101100000000000001011010110001111110001 :
(key == 10'b1000011111) ? 46'b1011010011100000000000001011010100000000111000 :
(key == 10'b1000100000) ? 46'b1011010001000000000000001011010001110010010010 :
(key == 10'b1000100001) ? 46'b1011001111000000000000001011001111100011111100 :
(key == 10'b1000100010) ? 46'b1011001101000000000000001011001101010101111000 :
(key == 10'b1000100011) ? 46'b1011001011000000000000001011001011001000000110 :
(key == 10'b1000100100) ? 46'b1011001000100000000000001011001000111010100101 :
(key == 10'b1000100101) ? 46'b1011000110000000000000001011000110101101010101 :
(key == 10'b1000100110) ? 46'b1011000100000000000000001011000100100000010110 :
(key == 10'b1000100111) ? 46'b1011000001100000000000001011000010010011101001 :
(key == 10'b1000101000) ? 46'b1010111111100000000000001011000000000111001100 :
(key == 10'b1000101001) ? 46'b1010111101100000000000001010111101111011000001 :
(key == 10'b1000101010) ? 46'b1010111011000000000000001010111011101111000111 :
(key == 10'b1000101011) ? 46'b1010111001000000000000001010111001100011011110 :
(key == 10'b1000101100) ? 46'b1010110111000000000000001010110111011000000101 :
(key == 10'b1000101101) ? 46'b1010110101000000000000001010110101001100111110 :
(key == 10'b1000101110) ? 46'b1010110010000000000000001010110011000010001000 :
(key == 10'b1000101111) ? 46'b1010110000000000000000001010110000110111100010 :
(key == 10'b1000110000) ? 46'b1010101110000000000000001010101110101101001101 :
(key == 10'b1000110001) ? 46'b1010101100000000000000001010101100100011001001 :
(key == 10'b1000110010) ? 46'b1010101010000000000000001010101010011001010101 :
(key == 10'b1000110011) ? 46'b1010100111100000000000001010101000001111110011 :
(key == 10'b1000110100) ? 46'b1010100110000000000000001010100110000110100000 :
(key == 10'b1000110101) ? 46'b1010100011100000000000001010100011111101011111 :
(key == 10'b1000110110) ? 46'b1010100001000000000000001010100001110100101110 :
(key == 10'b1000110111) ? 46'b1010011111100000000000001010011111101100001101 :
(key == 10'b1000111000) ? 46'b1010011101000000000000001010011101100011111101 :
(key == 10'b1000111001) ? 46'b1010011011000000000000001010011011011011111101 :
(key == 10'b1000111010) ? 46'b1010011001000000000000001010011001010100001110 :
(key == 10'b1000111011) ? 46'b1010010111000000000000001010010111001100101111 :
(key == 10'b1000111100) ? 46'b1010010100100000000000001010010101000101100001 :
(key == 10'b1000111101) ? 46'b1010010010100000000000001010010010111110100010 :
(key == 10'b1000111110) ? 46'b1010010000100000000000001010010000110111110100 :
(key == 10'b1000111111) ? 46'b1010001110100000000000001010001110110001010110 :
(key == 10'b1001000000) ? 46'b1010001100000000000000001010001100101011001000 :
(key == 10'b1001000001) ? 46'b1010001010100000000000001010001010100101001001 :
(key == 10'b1001000010) ? 46'b1010001000000000000000001010001000011111011100 :
(key == 10'b1001000011) ? 46'b1010000110100000000000001010000110011001111110 :
(key == 10'b1001000100) ? 46'b1010000100000000000000001010000100010100110001 :
(key == 10'b1001000101) ? 46'b1010000001100000000000001010000010001111110011 :
(key == 10'b1001000110) ? 46'b1001111111100000000000001010000000001011000101 :
(key == 10'b1001000111) ? 46'b1001111110000000000000001001111110000110100110 :
(key == 10'b1001001000) ? 46'b1001111011100000000000001001111100000010011000 :
(key == 10'b1001001001) ? 46'b1001111001100000000000001001111001111110011001 :
(key == 10'b1001001010) ? 46'b1001110111100000000000001001110111111010101010 :
(key == 10'b1001001011) ? 46'b1001110101100000000000001001110101110111001100 :
(key == 10'b1001001100) ? 46'b1001110011100000000000001001110011110011111011 :
(key == 10'b1001001101) ? 46'b1001110001100000000000001001110001110000111100 :
(key == 10'b1001001110) ? 46'b1001101111100000000000001001101111101110001011 :
(key == 10'b1001001111) ? 46'b1001101101000000000000001001101101101011101011 :
(key == 10'b1001010000) ? 46'b1001101011000000000000001001101011101001011010 :
(key == 10'b1001010001) ? 46'b1001101001000000000000001001101001100111010111 :
(key == 10'b1001010010) ? 46'b1001100111000000000000001001100111100101100101 :
(key == 10'b1001010011) ? 46'b1001100101000000000000001001100101100100000011 :
(key == 10'b1001010100) ? 46'b1001100011100000000000001001100011100010101110 :
(key == 10'b1001010101) ? 46'b1001100001000000000000001001100001100001101010 :
(key == 10'b1001010110) ? 46'b1001011111000000000000001001011111100000110101 :
(key == 10'b1001010111) ? 46'b1001011101000000000000001001011101100000001111 :
(key == 10'b1001011000) ? 46'b1001011011000000000000001001011011011111111000 :
(key == 10'b1001011001) ? 46'b1001011001000000000000001001011001011111110001 :
(key == 10'b1001011010) ? 46'b1001010111000000000000001001010111011111111000 :
(key == 10'b1001011011) ? 46'b1001010101000000000000001001010101100000001111 :
(key == 10'b1001011100) ? 46'b1001010011000000000000001001010011100000110100 :
(key == 10'b1001011101) ? 46'b1001010001000000000000001001010001100001101001 :
(key == 10'b1001011110) ? 46'b1001001111000000000000001001001111100010101101 :
(key == 10'b1001011111) ? 46'b1001001101000000000000001001001101100100000000 :
(key == 10'b1001100000) ? 46'b1001001011100000000000001001001011100101100001 :
(key == 10'b1001100001) ? 46'b1001001001000000000000001001001001100111010001 :
(key == 10'b1001100010) ? 46'b1001000111000000000000001001000111101001010001 :
(key == 10'b1001100011) ? 46'b1001000101000000000000001001000101101011011111 :
(key == 10'b1001100100) ? 46'b1001000011100000000000001001000011101101111011 :
(key == 10'b1001100101) ? 46'b1001000001000000000000001001000001110000100111 :
(key == 10'b1001100110) ? 46'b1000111111100000000000001000111111110011100001 :
(key == 10'b1001100111) ? 46'b1000111101100000000000001000111101110110101010 :
(key == 10'b1001101000) ? 46'b1000111011100000000000001000111011111010000001 :
(key == 10'b1001101001) ? 46'b1000111001100000000000001000111001111101100111 :
(key == 10'b1001101010) ? 46'b1000110111100000000000001000111000000001011011 :
(key == 10'b1001101011) ? 46'b1000110101100000000000001000110110000101011110 :
(key == 10'b1001101100) ? 46'b1000110011100000000000001000110100001001110000 :
(key == 10'b1001101101) ? 46'b1000110001100000000000001000110010001110010000 :
(key == 10'b1001101110) ? 46'b1000101111100000000000001000110000010010111110 :
(key == 10'b1001101111) ? 46'b1000101110000000000000001000101110010111111011 :
(key == 10'b1001110000) ? 46'b1000101100000000000000001000101100011101000110 :
(key == 10'b1001110001) ? 46'b1000101010000000000000001000101010100010011111 :
(key == 10'b1001110010) ? 46'b1000101000000000000000001000101000101000000111 :
(key == 10'b1001110011) ? 46'b1000100110100000000000001000100110101101111101 :
(key == 10'b1001110100) ? 46'b1000100100100000000000001000100100110100000001 :
(key == 10'b1001110101) ? 46'b1000100010100000000000001000100010111010010010 :
(key == 10'b1001110110) ? 46'b1000100000100000000000001000100001000000110011 :
(key == 10'b1001110111) ? 46'b1000011111000000000000001000011111000111100001 :
(key == 10'b1001111000) ? 46'b1000011100100000000000001000011101001110011110 :
(key == 10'b1001111001) ? 46'b1000011010100000000000001000011011010101101000 :
(key == 10'b1001111010) ? 46'b1000011001000000000000001000011001011101000000 :
(key == 10'b1001111011) ? 46'b1000010111000000000000001000010111100100100111 :
(key == 10'b1001111100) ? 46'b1000010101100000000000001000010101101100011010 :
(key == 10'b1001111101) ? 46'b1000010011100000000000001000010011110100011101 :
(key == 10'b1001111110) ? 46'b1000010001100000000000001000010001111100101101 :
(key == 10'b1001111111) ? 46'b1000001111100000000000001000010000000101001011 :
(key == 10'b1010000000) ? 46'b1000001101100000000000001000001110001101110110 :
(key == 10'b1010000001) ? 46'b1000001100000000000000001000001100010110110000 :
(key == 10'b1010000010) ? 46'b1000001010100000000000001000001010011111110110 :
(key == 10'b1010000011) ? 46'b1000001000000000000000001000001000101001001011 :
(key == 10'b1010000100) ? 46'b1000000110100000000000001000000110110010101110 :
(key == 10'b1010000101) ? 46'b1000000100100000000000001000000100111100011110 :
(key == 10'b1010000110) ? 46'b1000000010100000000000001000000011000110011100 :
(key == 10'b1010000111) ? 46'b1000000001000000000000001000000001010000100111 :
(key == 10'b1010001000) ? 46'b0111111110100000000000000111111111011011000000 :
(key == 10'b1010001001) ? 46'b0111111101000000000000000111111101100101100110 :
(key == 10'b1010001010) ? 46'b0111111011100000000000000111111011110000011001 :
(key == 10'b1010001011) ? 46'b0111111001100000000000000111111001111011011001 :
(key == 10'b1010001100) ? 46'b0111111000000000000000000111111000000110101000 :
(key == 10'b1010001101) ? 46'b0111110110000000000000000111110110010010000101 :
(key == 10'b1010001110) ? 46'b0111110100000000000000000111110100011101101101 :
(key == 10'b1010001111) ? 46'b0111110010000000000000000111110010101001100100 :
(key == 10'b1010010000) ? 46'b0111110000100000000000000111110000110101101000 :
(key == 10'b1010010001) ? 46'b0111101111000000000000000111101111000001111000 :
(key == 10'b1010010010) ? 46'b0111101100100000000000000111101101001110010111 :
(key == 10'b1010010011) ? 46'b0111101011000000000000000111101011011011000001 :
(key == 10'b1010010100) ? 46'b0111101001100000000000000111101001100111111010 :
(key == 10'b1010010101) ? 46'b0111100111100000000000000111100111110100111111 :
(key == 10'b1010010110) ? 46'b0111100101100000000000000111100110000010010011 :
(key == 10'b1010010111) ? 46'b0111100100000000000000000111100100001111110010 :
(key == 10'b1010011000) ? 46'b0111100010000000000000000111100010011101011111 :
(key == 10'b1010011001) ? 46'b0111100000100000000000000111100000101011011000 :
(key == 10'b1010011010) ? 46'b0111011110100000000000000111011110111001011111 :
(key == 10'b1010011011) ? 46'b0111011100100000000000000111011101000111110010 :
(key == 10'b1010011100) ? 46'b0111011011000000000000000111011011010110010011 :
(key == 10'b1010011101) ? 46'b0111011001100000000000000111011001100101000000 :
(key == 10'b1010011110) ? 46'b0111010111000000000000000111010111110011111011 :
(key == 10'b1010011111) ? 46'b0111010101100000000000000111010110000011000010 :
(key == 10'b1010100000) ? 46'b0111010100000000000000000111010100010010010101 :
(key == 10'b1010100001) ? 46'b0111010010000000000000000111010010100001110110 :
(key == 10'b1010100010) ? 46'b0111010000000000000000000111010000110001100011 :
(key == 10'b1010100011) ? 46'b0111001110100000000000000111001111000001011100 :
(key == 10'b1010100100) ? 46'b0111001100100000000000000111001101010001100011 :
(key == 10'b1010100101) ? 46'b0111001011000000000000000111001011100001110110 :
(key == 10'b1010100110) ? 46'b0111001001000000000000000111001001110010010111 :
(key == 10'b1010100111) ? 46'b0111000111100000000000000111001000000011000010 :
(key == 10'b1010101000) ? 46'b0111000110000000000000000111000110010011111011 :
(key == 10'b1010101001) ? 46'b0111000100100000000000000111000100100101000000 :
(key == 10'b1010101010) ? 46'b0111000010100000000000000111000010110110010011 :
(key == 10'b1010101011) ? 46'b0111000000100000000000000111000001000111110001 :
(key == 10'b1010101100) ? 46'b0110111111000000000000000110111111011001011100 :
(key == 10'b1010101101) ? 46'b0110111101100000000000000110111101101011010010 :
(key == 10'b1010101110) ? 46'b0110111011100000000000000110111011111101010110 :
(key == 10'b1010101111) ? 46'b0110111010000000000000000110111010001111100110 :
(key == 10'b1010110000) ? 46'b0110111000000000000000000110111000100010000001 :
(key == 10'b1010110001) ? 46'b0110110110000000000000000110110110110100101010 :
(key == 10'b1010110010) ? 46'b0110110100100000000000000110110101000111011111 :
(key == 10'b1010110011) ? 46'b0110110011000000000000000110110011011010100000 :
(key == 10'b1010110100) ? 46'b0110110001100000000000000110110001101101101100 :
(key == 10'b1010110101) ? 46'b0110101111100000000000000110110000000001000101 :
(key == 10'b1010110110) ? 46'b0110101110000000000000000110101110010100101010 :
(key == 10'b1010110111) ? 46'b0110101100100000000000000110101100101000011100 :
(key == 10'b1010111000) ? 46'b0110101010100000000000000110101010111100011001 :
(key == 10'b1010111001) ? 46'b0110101000100000000000000110101001010000100011 :
(key == 10'b1010111010) ? 46'b0110100111100000000000000110100111100100111000 :
(key == 10'b1010111011) ? 46'b0110100101100000000000000110100101111001011010 :
(key == 10'b1010111100) ? 46'b0110100100000000000000000110100100001110000111 :
(key == 10'b1010111101) ? 46'b0110100010100000000000000110100010100011000000 :
(key == 10'b1010111110) ? 46'b0110100000100000000000000110100000111000000111 :
(key == 10'b1010111111) ? 46'b0110011111000000000000000110011111001101010111 :
(key == 10'b1011000000) ? 46'b0110011101000000000000000110011101100010110100 :
(key == 10'b1011000001) ? 46'b0110011011100000000000000110011011111000011101 :
(key == 10'b1011000010) ? 46'b0110011010000000000000000110011010001110010010 :
(key == 10'b1011000011) ? 46'b0110011000100000000000000110011000100100010010 :
(key == 10'b1011000100) ? 46'b0110010110100000000000000110010110111010011110 :
(key == 10'b1011000101) ? 46'b0110010101000000000000000110010101010000110110 :
(key == 10'b1011000110) ? 46'b0110010011000000000000000110010011100111011010 :
(key == 10'b1011000111) ? 46'b0110010001100000000000000110010001111110001001 :
(key == 10'b1011001000) ? 46'b0110010000000000000000000110010000010101000011 :
(key == 10'b1011001001) ? 46'b0110001110100000000000000110001110101100001010 :
(key == 10'b1011001010) ? 46'b0110001100100000000000000110001101000011011101 :
(key == 10'b1011001011) ? 46'b0110001011000000000000000110001011011010111010 :
(key == 10'b1011001100) ? 46'b0110001001100000000000000110001001110010100011 :
(key == 10'b1011001101) ? 46'b0110000111100000000000000110001000001010011000 :
(key == 10'b1011001110) ? 46'b0110000110000000000000000110000110100010011000 :
(key == 10'b1011001111) ? 46'b0110000100100000000000000110000100111010100011 :
(key == 10'b1011010000) ? 46'b0110000011000000000000000110000011010010111011 :
(key == 10'b1011010001) ? 46'b0110000001000000000000000110000001101011011101 :
(key == 10'b1011010010) ? 46'b0101111111100000000000000110000000000100001010 :
(key == 10'b1011010011) ? 46'b0101111110100000000000000101111110011101000011 :
(key == 10'b1011010100) ? 46'b0101111100100000000000000101111100110110001000 :
(key == 10'b1011010101) ? 46'b0101111010100000000000000101111011001111011000 :
(key == 10'b1011010110) ? 46'b0101111001000000000000000101111001101000110011 :
(key == 10'b1011010111) ? 46'b0101111000000000000000000101111000000010011001 :
(key == 10'b1011011000) ? 46'b0101110101100000000000000101110110011100001011 :
(key == 10'b1011011001) ? 46'b0101110100100000000000000101110100110110000111 :
(key == 10'b1011011010) ? 46'b0101110010100000000000000101110011010000001111 :
(key == 10'b1011011011) ? 46'b0101110001000000000000000101110001101010100010 :
(key == 10'b1011011100) ? 46'b0101110000000000000000000101110000000100111111 :
(key == 10'b1011011101) ? 46'b0101101110000000000000000101101110011111101001 :
(key == 10'b1011011110) ? 46'b0101101101000000000000000101101100111010011101 :
(key == 10'b1011011111) ? 46'b0101101011000000000000000101101011010101011101 :
(key == 10'b1011100000) ? 46'b0101101001000000000000000101101001110000100111 :
(key == 10'b1011100001) ? 46'b0101101000000000000000000101101000001011111100 :
(key == 10'b1011100010) ? 46'b0101100110100000000000000101100110100111011100 :
(key == 10'b1011100011) ? 46'b0101100100100000000000000101100101000011000111 :
(key == 10'b1011100100) ? 46'b0101100011000000000000000101100011011110111110 :
(key == 10'b1011100101) ? 46'b0101100001100000000000000101100001111010111110 :
(key == 10'b1011100110) ? 46'b0101100000000000000000000101100000010111001011 :
(key == 10'b1011100111) ? 46'b0101011110100000000000000101011110110011100001 :
(key == 10'b1011101000) ? 46'b0101011101000000000000000101011101010000000010 :
(key == 10'b1011101001) ? 46'b0101011011100000000000000101011011101100101110 :
(key == 10'b1011101010) ? 46'b0101011010000000000000000101011010001001100101 :
(key == 10'b1011101011) ? 46'b0101011000000000000000000101011000100110100111 :
(key == 10'b1011101100) ? 46'b0101010110100000000000000101010111000011110100 :
(key == 10'b1011101101) ? 46'b0101010101000000000000000101010101100001001010 :
(key == 10'b1011101110) ? 46'b0101010100000000000000000101010011111110101100 :
(key == 10'b1011101111) ? 46'b0101010010000000000000000101010010011100011010 :
(key == 10'b1011110000) ? 46'b0101010000100000000000000101010000111010010000 :
(key == 10'b1011110001) ? 46'b0101001111100000000000000101001111011000010010 :
(key == 10'b1011110010) ? 46'b0101001101100000000000000101001101110110011111 :
(key == 10'b1011110011) ? 46'b0101001011100000000000000101001100010100110110 :
(key == 10'b1011110100) ? 46'b0101001010100000000000000101001010110011010110 :
(key == 10'b1011110101) ? 46'b0101001001000000000000000101001001010010000010 :
(key == 10'b1011110110) ? 46'b0101000111100000000000000101000111110000111001 :
(key == 10'b1011110111) ? 46'b0101000110000000000000000101000110001111111010 :
(key == 10'b1011111000) ? 46'b0101000100100000000000000101000100101111000101 :
(key == 10'b1011111001) ? 46'b0101000011000000000000000101000011001110011010 :
(key == 10'b1011111010) ? 46'b0101000001100000000000000101000001101101111010 :
(key == 10'b1011111011) ? 46'b0101000000000000000000000101000000001101100100 :
(key == 10'b1011111100) ? 46'b0100111110000000000000000100111110101101011010 :
(key == 10'b1011111101) ? 46'b0100111100100000000000000100111101001101011001 :
(key == 10'b1011111110) ? 46'b0100111011100000000000000100111011101101100010 :
(key == 10'b1011111111) ? 46'b0100111010000000000000000100111010001101110110 :
(key == 10'b1100000000) ? 46'b0100111000100000000000000100111000101110010011 :
(key == 10'b1100000001) ? 46'b0100110111000000000000000100110111001110111011 :
(key == 10'b1100000010) ? 46'b0100110101100000000000000100110101101111101101 :
(key == 10'b1100000011) ? 46'b0100110100000000000000000100110100010000101010 :
(key == 10'b1100000100) ? 46'b0100110010100000000000000100110010110001110001 :
(key == 10'b1100000101) ? 46'b0100110001000000000000000100110001010011000010 :
(key == 10'b1100000110) ? 46'b0100101111100000000000000100101111110100011101 :
(key == 10'b1100000111) ? 46'b0100101110000000000000000100101110010110000001 :
(key == 10'b1100001000) ? 46'b0100101100100000000000000100101100110111110000 :
(key == 10'b1100001001) ? 46'b0100101011100000000000000100101011011001101001 :
(key == 10'b1100001010) ? 46'b0100101001100000000000000100101001111011101101 :
(key == 10'b1100001011) ? 46'b0100101000000000000000000100101000011101111010 :
(key == 10'b1100001100) ? 46'b0100100111000000000000000100100111000000010001 :
(key == 10'b1100001101) ? 46'b0100100101000000000000000100100101100010110010 :
(key == 10'b1100001110) ? 46'b0100100011100000000000000100100100000101011101 :
(key == 10'b1100001111) ? 46'b0100100010100000000000000100100010101000010001 :
(key == 10'b1100010000) ? 46'b0100100001000000000000000100100001001011010001 :
(key == 10'b1100010001) ? 46'b0100011111000000000000000100011111101110011001 :
(key == 10'b1100010010) ? 46'b0100011110000000000000000100011110010001101011 :
(key == 10'b1100010011) ? 46'b0100011100100000000000000100011100110101001000 :
(key == 10'b1100010100) ? 46'b0100011011000000000000000100011011011000101101 :
(key == 10'b1100010101) ? 46'b0100011001100000000000000100011001111100011110 :
(key == 10'b1100010110) ? 46'b0100011000000000000000000100011000100000010111 :
(key == 10'b1100010111) ? 46'b0100010110100000000000000100010111000100011011 :
(key == 10'b1100011000) ? 46'b0100010101100000000000000100010101101000100111 :
(key == 10'b1100011001) ? 46'b0100010100000000000000000100010100001100111110 :
(key == 10'b1100011010) ? 46'b0100010011000000000000000100010010110001011110 :
(key == 10'b1100011011) ? 46'b0100010001000000000000000100010001010110001001 :
(key == 10'b1100011100) ? 46'b0100001111100000000000000100001111111010111101 :
(key == 10'b1100011101) ? 46'b0100001110000000000000000100001110011111111010 :
(key == 10'b1100011110) ? 46'b0100001100100000000000000100001101000101000001 :
(key == 10'b1100011111) ? 46'b0100001011100000000000000100001011101010010001 :
(key == 10'b1100100000) ? 46'b0100001010000000000000000100001010001111101011 :
(key == 10'b1100100001) ? 46'b0100001000100000000000000100001000110101001111 :
(key == 10'b1100100010) ? 46'b0100000111000000000000000100000111011010111100 :
(key == 10'b1100100011) ? 46'b0100000101100000000000000100000110000000110011 :
(key == 10'b1100100100) ? 46'b0100000100000000000000000100000100100110110011 :
(key == 10'b1100100101) ? 46'b0100000011000000000000000100000011001100111100 :
(key == 10'b1100100110) ? 46'b0100000001100000000000000100000001110011001111 :
(key == 10'b1100100111) ? 46'b0100000000000000000000000100000000011001101100 :
(key == 10'b1100101000) ? 46'b0011111110100000000000000011111111000000010001 :
(key == 10'b1100101001) ? 46'b0011111101000000000000000011111101100111000000 :
(key == 10'b1100101010) ? 46'b0011111011100000000000000011111100001101111000 :
(key == 10'b1100101011) ? 46'b0011111010100000000000000011111010110100111010 :
(key == 10'b1100101100) ? 46'b0011111001000000000000000011111001011100000100 :
(key == 10'b1100101101) ? 46'b0011111000000000000000000011111000000011011001 :
(key == 10'b1100101110) ? 46'b0011110110000000000000000011110110101010110111 :
(key == 10'b1100101111) ? 46'b0011110101000000000000000011110101010010011101 :
(key == 10'b1100110000) ? 46'b0011110011100000000000000011110011111010001110 :
(key == 10'b1100110001) ? 46'b0011110010000000000000000011110010100010000111 :
(key == 10'b1100110010) ? 46'b0011110001000000000000000011110001001010001001 :
(key == 10'b1100110011) ? 46'b0011101111100000000000000011101111110010010100 :
(key == 10'b1100110100) ? 46'b0011101110000000000000000011101110011010101001 :
(key == 10'b1100110101) ? 46'b0011101100100000000000000011101101000011000111 :
(key == 10'b1100110110) ? 46'b0011101011000000000000000011101011101011101110 :
(key == 10'b1100110111) ? 46'b0011101010000000000000000011101010010100011110 :
(key == 10'b1100111000) ? 46'b0011101000100000000000000011101000111101010111 :
(key == 10'b1100111001) ? 46'b0011100111000000000000000011100111100110011001 :
(key == 10'b1100111010) ? 46'b0011100110000000000000000011100110001111100011 :
(key == 10'b1100111011) ? 46'b0011100100100000000000000011100100111000111000 :
(key == 10'b1100111100) ? 46'b0011100011000000000000000011100011100010010101 :
(key == 10'b1100111101) ? 46'b0011100001100000000000000011100010001011111011 :
(key == 10'b1100111110) ? 46'b0011100000100000000000000011100000110101101010 :
(key == 10'b1100111111) ? 46'b0011011111000000000000000011011111011111100010 :
(key == 10'b1101000000) ? 46'b0011011101100000000000000011011110001001100011 :
(key == 10'b1101000001) ? 46'b0011011100100000000000000011011100110011101100 :
(key == 10'b1101000010) ? 46'b0011011011100000000000000011011011011101111110 :
(key == 10'b1101000011) ? 46'b0011011010000000000000000011011010001000011010 :
(key == 10'b1101000100) ? 46'b0011011000100000000000000011011000110010111110 :
(key == 10'b1101000101) ? 46'b0011010111000000000000000011010111011101101100 :
(key == 10'b1101000110) ? 46'b0011010101100000000000000011010110001000100010 :
(key == 10'b1101000111) ? 46'b0011010100100000000000000011010100110011100000 :
(key == 10'b1101001000) ? 46'b0011010011000000000000000011010011011110100111 :
(key == 10'b1101001001) ? 46'b0011010001100000000000000011010010001001110111 :
(key == 10'b1101001010) ? 46'b0011010000100000000000000011010000110101010000 :
(key == 10'b1101001011) ? 46'b0011001111100000000000000011001111100000110001 :
(key == 10'b1101001100) ? 46'b0011001110000000000000000011001110001100011100 :
(key == 10'b1101001101) ? 46'b0011001100100000000000000011001100111000001111 :
(key == 10'b1101001110) ? 46'b0011001011000000000000000011001011100100001010 :
(key == 10'b1101001111) ? 46'b0011001010000000000000000011001010010000001110 :
(key == 10'b1101010000) ? 46'b0011001000100000000000000011001000111100011011 :
(key == 10'b1101010001) ? 46'b0011000111100000000000000011000111101000110000 :
(key == 10'b1101010010) ? 46'b0011000110000000000000000011000110010101001110 :
(key == 10'b1101010011) ? 46'b0011000100100000000000000011000101000001110100 :
(key == 10'b1101010100) ? 46'b0011000011100000000000000011000011101110100011 :
(key == 10'b1101010101) ? 46'b0011000010000000000000000011000010011011011011 :
(key == 10'b1101010110) ? 46'b0011000000100000000000000011000001001000011011 :
(key == 10'b1101010111) ? 46'b0010111111100000000000000010111111110101100011 :
(key == 10'b1101011000) ? 46'b0010111110100000000000000010111110100010110100 :
(key == 10'b1101011001) ? 46'b0010111101000000000000000010111101010000001110 :
(key == 10'b1101011010) ? 46'b0010111011100000000000000010111011111101101111 :
(key == 10'b1101011011) ? 46'b0010111010000000000000000010111010101011011001 :
(key == 10'b1101011100) ? 46'b0010111001000000000000000010111001011001001100 :
(key == 10'b1101011101) ? 46'b0010110111100000000000000010111000000111000111 :
(key == 10'b1101011110) ? 46'b0010110110100000000000000010110110110101001010 :
(key == 10'b1101011111) ? 46'b0010110101000000000000000010110101100011010101 :
(key == 10'b1101100000) ? 46'b0010110100100000000000000010110100010001101001 :
(key == 10'b1101100001) ? 46'b0010110010100000000000000010110011000000000110 :
(key == 10'b1101100010) ? 46'b0010110001100000000000000010110001101110101001 :
(key == 10'b1101100011) ? 46'b0010110000000000000000000010110000011101010111 :
(key == 10'b1101100100) ? 46'b0010101111000000000000000010101111001100001100 :
(key == 10'b1101100101) ? 46'b0010101101100000000000000010101101111011001001 :
(key == 10'b1101100110) ? 46'b0010101100100000000000000010101100101010001110 :
(key == 10'b1101100111) ? 46'b0010101011100000000000000010101011011001011100 :
(key == 10'b1101101000) ? 46'b0010101010000000000000000010101010001000110010 :
(key == 10'b1101101001) ? 46'b0010101000100000000000000010101000111000010000 :
(key == 10'b1101101010) ? 46'b0010100111100000000000000010100111100111110110 :
(key == 10'b1101101011) ? 46'b0010100110000000000000000010100110010111100100 :
(key == 10'b1101101100) ? 46'b0010100101000000000000000010100101000111011010 :
(key == 10'b1101101101) ? 46'b0010100011100000000000000010100011110111011001 :
(key == 10'b1101101110) ? 46'b0010100010100000000000000010100010100111011111 :
(key == 10'b1101101111) ? 46'b0010100001000000000000000010100001010111101110 :
(key == 10'b1101110000) ? 46'b0010100000000000000000000010100000001000000100 :
(key == 10'b1101110001) ? 46'b0010011111000000000000000010011110111000100011 :
(key == 10'b1101110010) ? 46'b0010011101100000000000000010011101101001001001 :
(key == 10'b1101110011) ? 46'b0010011100000000000000000010011100011001111000 :
(key == 10'b1101110100) ? 46'b0010011011000000000000000010011011001010101111 :
(key == 10'b1101110101) ? 46'b0010011001100000000000000010011001111011101110 :
(key == 10'b1101110110) ? 46'b0010011000000000000000000010011000101100110100 :
(key == 10'b1101110111) ? 46'b0010010111100000000000000010010111011110000010 :
(key == 10'b1101111000) ? 46'b0010010110000000000000000010010110001111011001 :
(key == 10'b1101111001) ? 46'b0010010101000000000000000010010101000000110111 :
(key == 10'b1101111010) ? 46'b0010010011100000000000000010010011110010011101 :
(key == 10'b1101111011) ? 46'b0010010010000000000000000010010010100100001011 :
(key == 10'b1101111100) ? 46'b0010010001000000000000000010010001010110000000 :
(key == 10'b1101111101) ? 46'b0010010000000000000000000010010000000111111110 :
(key == 10'b1101111110) ? 46'b0010001111000000000000000010001110111010000011 :
(key == 10'b1101111111) ? 46'b0010001101100000000000000010001101101100010001 :
(key == 10'b1110000000) ? 46'b0010001100000000000000000010001100011110100110 :
(key == 10'b1110000001) ? 46'b0010001011000000000000000010001011010001000010 :
(key == 10'b1110000010) ? 46'b0010001010000000000000000010001010000011100110 :
(key == 10'b1110000011) ? 46'b0010001000100000000000000010001000110110010100 :
(key == 10'b1110000100) ? 46'b0010000111000000000000000010000111101001000111 :
(key == 10'b1110000101) ? 46'b0010000110100000000000000010000110011100000010 :
(key == 10'b1110000110) ? 46'b0010000101000000000000000010000101001111000110 :
(key == 10'b1110000111) ? 46'b0010000011100000000000000010000100000010010001 :
(key == 10'b1110001000) ? 46'b0010000010100000000000000010000010110101100100 :
(key == 10'b1110001001) ? 46'b0010000001000000000000000010000001101000111110 :
(key == 10'b1110001010) ? 46'b0010000000000000000000000010000000011100100000 :
(key == 10'b1110001011) ? 46'b0001111111000000000000000001111111010000001001 :
(key == 10'b1110001100) ? 46'b0001111101100000000000000001111110000011111010 :
(key == 10'b1110001101) ? 46'b0001111100100000000000000001111100110111110011 :
(key == 10'b1110001110) ? 46'b0001111011100000000000000001111011101011110011 :
(key == 10'b1110001111) ? 46'b0001111010100000000000000001111010011111111010 :
(key == 10'b1110010000) ? 46'b0001111001000000000000000001111001010100001010 :
(key == 10'b1110010001) ? 46'b0001110111100000000000000001111000001000100001 :
(key == 10'b1110010010) ? 46'b0001110110100000000000000001110110111100111111 :
(key == 10'b1110010011) ? 46'b0001110101100000000000000001110101110001100100 :
(key == 10'b1110010100) ? 46'b0001110100100000000000000001110100100110010001 :
(key == 10'b1110010101) ? 46'b0001110011000000000000000001110011011011000101 :
(key == 10'b1110010110) ? 46'b0001110010000000000000000001110010010000000010 :
(key == 10'b1110010111) ? 46'b0001110001000000000000000001110001000101000101 :
(key == 10'b1110011000) ? 46'b0001110000000000000000000001101111111010010000 :
(key == 10'b1110011001) ? 46'b0001101110100000000000000001101110101111100010 :
(key == 10'b1110011010) ? 46'b0001101101000000000000000001101101100100111100 :
(key == 10'b1110011011) ? 46'b0001101100000000000000000001101100011010011101 :
(key == 10'b1110011100) ? 46'b0001101011000000000000000001101011010000000101 :
(key == 10'b1110011101) ? 46'b0001101001100000000000000001101010000101110101 :
(key == 10'b1110011110) ? 46'b0001101001000000000000000001101000111011101011 :
(key == 10'b1110011111) ? 46'b0001100111100000000000000001100111110001101010 :
(key == 10'b1110100000) ? 46'b0001100110100000000000000001100110100111101111 :
(key == 10'b1110100001) ? 46'b0001100101000000000000000001100101011101111100 :
(key == 10'b1110100010) ? 46'b0001100100000000000000000001100100010100010000 :
(key == 10'b1110100011) ? 46'b0001100010100000000000000001100011001010101100 :
(key == 10'b1110100100) ? 46'b0001100010000000000000000001100010000001001101 :
(key == 10'b1110100101) ? 46'b0001100001000000000000000001100000110111110111 :
(key == 10'b1110100110) ? 46'b0001011111100000000000000001011111101110101000 :
(key == 10'b1110100111) ? 46'b0001011110000000000000000001011110100101100001 :
(key == 10'b1110101000) ? 46'b0001011101100000000000000001011101011100011111 :
(key == 10'b1110101001) ? 46'b0001011100000000000000000001011100010011100101 :
(key == 10'b1110101010) ? 46'b0001011011000000000000000001011011001010110011 :
(key == 10'b1110101011) ? 46'b0001011001100000000000000001011010000010001000 :
(key == 10'b1110101100) ? 46'b0001011000100000000000000001011000111001100011 :
(key == 10'b1110101101) ? 46'b0001011000000000000000000001010111110001000101 :
(key == 10'b1110101110) ? 46'b0001010110000000000000000001010110101000110000 :
(key == 10'b1110101111) ? 46'b0001010101100000000000000001010101100000100000 :
(key == 10'b1110110000) ? 46'b0001010100000000000000000001010100011000011001 :
(key == 10'b1110110001) ? 46'b0001010011000000000000000001010011010000010111 :
(key == 10'b1110110010) ? 46'b0001010001100000000000000001010010001000011110 :
(key == 10'b1110110011) ? 46'b0001010001000000000000000001010001000000101010 :
(key == 10'b1110110100) ? 46'b0001010000000000000000000001001111111000111110 :
(key == 10'b1110110101) ? 46'b0001001110100000000000000001001110110001011001 :
(key == 10'b1110110110) ? 46'b0001001101100000000000000001001101101001111011 :
(key == 10'b1110110111) ? 46'b0001001100000000000000000001001100100010100100 :
(key == 10'b1110111000) ? 46'b0001001011000000000000000001001011011011010100 :
(key == 10'b1110111001) ? 46'b0001001010100000000000000001001010010100001010 :
(key == 10'b1110111010) ? 46'b0001001001000000000000000001001001001101000111 :
(key == 10'b1110111011) ? 46'b0001000111100000000000000001001000000110001100 :
(key == 10'b1110111100) ? 46'b0001000110100000000000000001000110111111011000 :
(key == 10'b1110111101) ? 46'b0001000101100000000000000001000101111000101010 :
(key == 10'b1110111110) ? 46'b0001000100000000000000000001000100110010000011 :
(key == 10'b1110111111) ? 46'b0001000011000000000000000001000011101011100011 :
(key == 10'b1111000000) ? 46'b0001000010100000000000000001000010100101001001 :
(key == 10'b1111000001) ? 46'b0001000001000000000000000001000001011110110111 :
(key == 10'b1111000010) ? 46'b0001000000000000000000000001000000011000101011 :
(key == 10'b1111000011) ? 46'b0000111111000000000000000000111111010010100110 :
(key == 10'b1111000100) ? 46'b0000111110000000000000000000111110001100101000 :
(key == 10'b1111000101) ? 46'b0000111101000000000000000000111101000110110000 :
(key == 10'b1111000110) ? 46'b0000111011100000000000000000111100000001000000 :
(key == 10'b1111000111) ? 46'b0000111010100000000000000000111010111011010110 :
(key == 10'b1111001000) ? 46'b0000111001100000000000000000111001110101110011 :
(key == 10'b1111001001) ? 46'b0000111001000000000000000000111000110000010110 :
(key == 10'b1111001010) ? 46'b0000110111000000000000000000110111101011000001 :
(key == 10'b1111001011) ? 46'b0000110110100000000000000000110110100101110001 :
(key == 10'b1111001100) ? 46'b0000110101000000000000000000110101100000101001 :
(key == 10'b1111001101) ? 46'b0000110100000000000000000000110100011011100111 :
(key == 10'b1111001110) ? 46'b0000110011000000000000000000110011010110101011 :
(key == 10'b1111001111) ? 46'b0000110010000000000000000000110010010001110111 :
(key == 10'b1111010000) ? 46'b0000110001000000000000000000110001001101001000 :
(key == 10'b1111010001) ? 46'b0000101111100000000000000000110000001000100010 :
(key == 10'b1111010010) ? 46'b0000101111000000000000000000101111000100000000 :
(key == 10'b1111010011) ? 46'b0000101101100000000000000000101101111111100110 :
(key == 10'b1111010100) ? 46'b0000101100100000000000000000101100111011010010 :
(key == 10'b1111010101) ? 46'b0000101011100000000000000000101011110111000101 :
(key == 10'b1111010110) ? 46'b0000101010100000000000000000101010110010111110 :
(key == 10'b1111010111) ? 46'b0000101001100000000000000000101001101110111110 :
(key == 10'b1111011000) ? 46'b0000101000100000000000000000101000101011000100 :
(key == 10'b1111011001) ? 46'b0000100111000000000000000000100111100111010001 :
(key == 10'b1111011010) ? 46'b0000100110100000000000000000100110100011100100 :
(key == 10'b1111011011) ? 46'b0000100101100000000000000000100101011111111110 :
(key == 10'b1111011100) ? 46'b0000100100100000000000000000100100011100011110 :
(key == 10'b1111011101) ? 46'b0000100011000000000000000000100011011001000101 :
(key == 10'b1111011110) ? 46'b0000100010100000000000000000100010010101110010 :
(key == 10'b1111011111) ? 46'b0000100001000000000000000000100001010010100101 :
(key == 10'b1111100000) ? 46'b0000100000000000000000000000100000001111011111 :
(key == 10'b1111100001) ? 46'b0000011111000000000000000000011111001100011111 :
(key == 10'b1111100010) ? 46'b0000011110000000000000000000011110001001100110 :
(key == 10'b1111100011) ? 46'b0000011101000000000000000000011101000110110011 :
(key == 10'b1111100100) ? 46'b0000011011100000000000000000011100000100000111 :
(key == 10'b1111100101) ? 46'b0000011011000000000000000000011011000001100000 :
(key == 10'b1111100110) ? 46'b0000011010000000000000000000011001111111000000 :
(key == 10'b1111100111) ? 46'b0000011000100000000000000000011000111100100111 :
(key == 10'b1111101000) ? 46'b0000010111100000000000000000010111111010010011 :
(key == 10'b1111101001) ? 46'b0000010110100000000000000000010110111000000101 :
(key == 10'b1111101010) ? 46'b0000010101100000000000000000010101110101111111 :
(key == 10'b1111101011) ? 46'b0000010100000000000000000000010100110011111111 :
(key == 10'b1111101100) ? 46'b0000010011100000000000000000010011110010000011 :
(key == 10'b1111101101) ? 46'b0000010010100000000000000000010010110000001111 :
(key == 10'b1111101110) ? 46'b0000010001100000000000000000010001101110100001 :
(key == 10'b1111101111) ? 46'b0000010000100000000000000000010000101100111001 :
(key == 10'b1111110000) ? 46'b0000001111100000000000000000001111101011011001 :
(key == 10'b1111110001) ? 46'b0000001110100000000000000000001110101001111101 :
(key == 10'b1111110010) ? 46'b0000001101100000000000000000001101101000100111 :
(key == 10'b1111110011) ? 46'b0000001100100000000000000000001100100111011001 :
(key == 10'b1111110100) ? 46'b0000001011000000000000000000001011100110010001 :
(key == 10'b1111110101) ? 46'b0000001010100000000000000000001010100101001101 :
(key == 10'b1111110110) ? 46'b0000001001100000000000000000001001100100010001 :
(key == 10'b1111110111) ? 46'b0000001000000000000000000000001000100011011011 :
(key == 10'b1111111000) ? 46'b0000000111100000000000000000000111100010101001 :
(key == 10'b1111111001) ? 46'b0000000110100000000000000000000110100001111111 :
(key == 10'b1111111010) ? 46'b0000000101100000000000000000000101100001011011 :
(key == 10'b1111111011) ? 46'b0000000100100000000000000000000100100000111101 :
(key == 10'b1111111100) ? 46'b0000000011100000000000000000000011100000100101 :
(key == 10'b1111111101) ? 46'b0000000010100000000000000000000010100000010011 :
(key == 10'b1111111110) ? 46'b0000000001100000000000000000000001100000000111 :
(key == 10'b1111111111) ? 46'b0000000000100000000000000000000000100000000001 : 46'd0;

endmodule

`default_nettype wire
