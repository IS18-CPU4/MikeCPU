`default_nettype none

module fsqrt_p2
   ( input wire [31:0] x,
     output reg [31:0] y,
     input wire clk,
     input wire rstn);

   // split sequence to each subsequence
   wire xs;
   wire [7:0] xe;
   wire [22:0] xm;
   reg [7:0] xe_r;
   reg [22:0] xm_r;
   assign {xs, xe, xm} = x;

   wire [7:0] shift_xe;
   assign shift_xe = xe >> 1;

   // calc e
   wire [7:0] e;
   reg [7:0] e_r;
   assign e = (xe[0] == 1) ? 8'd189 - shift_xe : 8'd190 - shift_xe; 

   // calc m
   wire [47:0] val;
   wire [10:0] key;
   assign key = {xe[0], xm[22:13]};

   // lookup table and get constant and grad
   lookup_table lt(key, val);


   wire [24:0] constant;
   reg [24:0] constant_r;
   wire [22:0] grad;
   assign constant = val[47:23];
   assign grad = val[22:0];

   wire [47:0] grad2;
   reg [47:0] grad2_r;
   assign grad2 = {1'b1, grad} * {1'b1, xm};

   // register insertion here
   
   wire [24:0] grad3_even;
   assign grad3_even = (grad2_r[47] == 1'b1) ? {2'd0, grad2_r[47:25]} :
                       (xm_r[22:13] != 10'b1111111111) ? {2'd0, grad2_r[46:24]} : {2'd0, grad2_r[47:25]};

   wire [24:0] grad3_odd;
   assign grad3_odd = (grad2_r[47] == 1'b0) ? {2'd0, grad2_r[46:24]} :
                      (xm_r[22:13] != 10'd0) ? {2'd0, grad2_r[47:25]} : {2'd0, grad2_r[46:24]};

   wire [24:0] tmp_m;
   assign tmp_m = (xe_r[0] == 1) ? constant_r - grad3_odd : constant_r - grad3_even;

   wire [22:0] m;
   assign m = tmp_m[22:0]; // ignore implicit 1

   wire [31:0] y_w;
   wire ovf;
   fmul u1({1'b0, xe_r, xm_r}, {1'b0, e_r, m}, y_w, ovf); // sign is 0

   always @(posedge clk) begin
    if (~rstn) begin
      y <= 0;
      xe_r <= 0;
      xm_r <= 0;
      e_r <= 0;
      constant_r <= 0;
      grad2_r <= 0;
    end else begin
      y <= y_w;
      xe_r <= xe;
      xm_r <= xm;
      e_r <= e;
      constant_r <= constant;
      grad2_r <= grad2;
    end
   end

endmodule

module lookup_table
   ( input wire [10:0] key,
     output wire [47:0] value);

   assign value =
(key == 11'b00000000000) ? 48'b100001111011101100111100001101001110001100001011 :
(key == 11'b00000000001) ? 48'b100001111010101001001010001101001001111101010100 :
(key == 11'b00000000010) ? 48'b100001111001100101011110001101000101101111000101 :
(key == 11'b00000000011) ? 48'b100001111000100001111000001101000001100001100011 :
(key == 11'b00000000100) ? 48'b100001110111011110011010001100111101010100101100 :
(key == 11'b00000000101) ? 48'b100001110110011011000001001100111001001000011011 :
(key == 11'b00000000110) ? 48'b100001110101010111101110001100110100111100110101 :
(key == 11'b00000000111) ? 48'b100001110100010100100010001100110000110001111011 :
(key == 11'b00000001000) ? 48'b100001110011010001011100001100101100100111100110 :
(key == 11'b00000001001) ? 48'b100001110010001110011100001100101000011101111101 :
(key == 11'b00000001010) ? 48'b100001110001001011100010001100100100010100111011 :
(key == 11'b00000001011) ? 48'b100001110000001000101111001100100000001100100010 :
(key == 11'b00000001100) ? 48'b100001101111000110000010001100011100000100110100 :
(key == 11'b00000001101) ? 48'b100001101110000011011100001100010111111101110000 :
(key == 11'b00000001110) ? 48'b100001101101000000111010001100010011110111001111 :
(key == 11'b00000001111) ? 48'b100001101011111110011111001100001111110001011001 :
(key == 11'b00000010000) ? 48'b100001101010111100001010001100001011101100001101 :
(key == 11'b00000010001) ? 48'b100001101001111001111100001100000111100111101001 :
(key == 11'b00000010010) ? 48'b100001101000110111110100001100000011100011101100 :
(key == 11'b00000010011) ? 48'b100001100111110101110010001011111111100000010111 :
(key == 11'b00000010100) ? 48'b100001100110110011110110001011111011011101101010 :
(key == 11'b00000010101) ? 48'b100001100101110001111111001011110111011011100011 :
(key == 11'b00000010110) ? 48'b100001100100110000001110001011110011011010000010 :
(key == 11'b00000010111) ? 48'b100001100011101110100100001011101111011001001010 :
(key == 11'b00000011000) ? 48'b100001100010101101000000001011101011011000111100 :
(key == 11'b00000011001) ? 48'b100001100001101011100011001011100111011001010101 :
(key == 11'b00000011010) ? 48'b100001100000101010001011001011100011011010010010 :
(key == 11'b00000011011) ? 48'b100001011111101000111000001011011111011011110111 :
(key == 11'b00000011100) ? 48'b100001011110100111101100001011011011011101111111 :
(key == 11'b00000011101) ? 48'b100001011101100110100101001011010111100000110001 :
(key == 11'b00000011110) ? 48'b100001011100100101100110001011010011100100001101 :
(key == 11'b00000011111) ? 48'b100001011011100100101011001011001111101000001010 :
(key == 11'b00000100000) ? 48'b100001011010100011110110001011001011101100101111 :
(key == 11'b00000100001) ? 48'b100001011001100011001000001011000111110001111000 :
(key == 11'b00000100010) ? 48'b100001011000100010011111001011000011110111101011 :
(key == 11'b00000100011) ? 48'b100001010111100001111101001010111111111110000100 :
(key == 11'b00000100100) ? 48'b100001010110100001100000001010111100000101000000 :
(key == 11'b00000100101) ? 48'b100001010101100001001000001010111000001100100000 :
(key == 11'b00000100110) ? 48'b100001010100100000110111001010110100010100101001 :
(key == 11'b00000100111) ? 48'b100001010011100000101100001010110000011101010100 :
(key == 11'b00000101000) ? 48'b100001010010100000100101001010101100100110100100 :
(key == 11'b00000101001) ? 48'b100001010001100000100101001010101000110000011011 :
(key == 11'b00000101010) ? 48'b100001010000100000101011001010100100111010110110 :
(key == 11'b00000101011) ? 48'b100001001111100000110110001010100001000101110110 :
(key == 11'b00000101100) ? 48'b100001001110100001001000001010011101010001011100 :
(key == 11'b00000101101) ? 48'b100001001101100001011110001010011001011101100110 :
(key == 11'b00000101110) ? 48'b100001001100100001111100001010010101101010010111 :
(key == 11'b00000101111) ? 48'b100001001011100010011110001010010001110111101000 :
(key == 11'b00000110000) ? 48'b100001001010100011000110001010001110000101011110 :
(key == 11'b00000110001) ? 48'b100001001001100011110011001010001010010011110111 :
(key == 11'b00000110010) ? 48'b100001001000100100100111001010000110100010111000 :
(key == 11'b00000110011) ? 48'b100001000111100101100000001010000010110010011000 :
(key == 11'b00000110100) ? 48'b100001000110100110011110001001111111000010011110 :
(key == 11'b00000110101) ? 48'b100001000101100111100011001001111011010011001001 :
(key == 11'b00000110110) ? 48'b100001000100101000101101001001110111100100011001 :
(key == 11'b00000110111) ? 48'b100001000011101001111100001001110011110110000101 :
(key == 11'b00000111000) ? 48'b100001000010101011010000001001110000001000011001 :
(key == 11'b00000111001) ? 48'b100001000001101100101100001001101100011011010010 :
(key == 11'b00000111010) ? 48'b100001000000101110001100001001101000101110101100 :
(key == 11'b00000111011) ? 48'b100000111111101111110001001001100101000010101000 :
(key == 11'b00000111100) ? 48'b100000111110110001011101001001100001010111001010 :
(key == 11'b00000111101) ? 48'b100000111101110011001110001001011101101100001100 :
(key == 11'b00000111110) ? 48'b100000111100110101000100001001011010000001110001 :
(key == 11'b00000111111) ? 48'b100000111011110111000000001001010110010111111010 :
(key == 11'b00001000000) ? 48'b100000111010111001000001001001010010101110100100 :
(key == 11'b00001000001) ? 48'b100000111001111011000111001001001111000101110000 :
(key == 11'b00001000010) ? 48'b100000111000111101010011001001001011011101011101 :
(key == 11'b00001000011) ? 48'b100000110111111111100110001001000111110101110001 :
(key == 11'b00001000100) ? 48'b100000110111000001111100001001000100001110100001 :
(key == 11'b00001000101) ? 48'b100000110110000100011000001001000000100111110101 :
(key == 11'b00001000110) ? 48'b100000110101000110111010001000111101000001101010 :
(key == 11'b00001000111) ? 48'b100000110100001001100001001000111001011100000011 :
(key == 11'b00001001000) ? 48'b100000110011001100001101001000110101110110111010 :
(key == 11'b00001001001) ? 48'b100000110010001111000000001000110010010010011000 :
(key == 11'b00001001010) ? 48'b100000110001010001110111001000101110101110010100 :
(key == 11'b00001001011) ? 48'b100000110000010100110011001000101011001010101101 :
(key == 11'b00001001100) ? 48'b100000101111010111110100001000100111100111101011 :
(key == 11'b00001001101) ? 48'b100000101110011010111100001000100100000101001100 :
(key == 11'b00001001110) ? 48'b100000101101011110001001001000100000100011001101 :
(key == 11'b00001001111) ? 48'b100000101100100001011011001000011101000001101101 :
(key == 11'b00001010000) ? 48'b100000101011100100110010001000011001100000101111 :
(key == 11'b00001010001) ? 48'b100000101010101000001110001000010110000000010000 :
(key == 11'b00001010010) ? 48'b100000101001101011110000001000010010100000010100 :
(key == 11'b00001010011) ? 48'b100000101000101111010111001000001111000000110101 :
(key == 11'b00001010100) ? 48'b100000100111110011000011001000001011100001111001 :
(key == 11'b00001010101) ? 48'b100000100110110110110100001000001000000011011011 :
(key == 11'b00001010110) ? 48'b100000100101111010101010001000000100100101011110 :
(key == 11'b00001010111) ? 48'b100000100100111110100111001000000001001000000010 :
(key == 11'b00001011000) ? 48'b100000100100000010101000000111111101101011000100 :
(key == 11'b00001011001) ? 48'b100000100011000110101101000111111010001110100100 :
(key == 11'b00001011010) ? 48'b100000100010001010111000000111110110110010100110 :
(key == 11'b00001011011) ? 48'b100000100001001111001001000111110011010111001011 :
(key == 11'b00001011100) ? 48'b100000100000010011011110000111101111111100001011 :
(key == 11'b00001011101) ? 48'b100000011111010111111001000111101100100001101100 :
(key == 11'b00001011110) ? 48'b100000011110011100011001000111101001000111101100 :
(key == 11'b00001011111) ? 48'b100000011101100000111110000111100101101110001010 :
(key == 11'b00001100000) ? 48'b100000011100100101101000000111100010010101001000 :
(key == 11'b00001100001) ? 48'b100000011011101010010111000111011110111100100110 :
(key == 11'b00001100010) ? 48'b100000011010101111001011000111011011100100100011 :
(key == 11'b00001100011) ? 48'b100000011001110100000100000111011000001100111101 :
(key == 11'b00001100100) ? 48'b100000011000111001000010000111010100110101110110 :
(key == 11'b00001100101) ? 48'b100000010111111110000110000111010001011111001111 :
(key == 11'b00001100110) ? 48'b100000010111000011001110000111001110001001000101 :
(key == 11'b00001100111) ? 48'b100000010110001000011011000111001010110011011001 :
(key == 11'b00001101000) ? 48'b100000010101001101101101000111000111011110001010 :
(key == 11'b00001101001) ? 48'b100000010100010011000101000111000100001001011101 :
(key == 11'b00001101010) ? 48'b100000010011011000100001000111000000110101001100 :
(key == 11'b00001101011) ? 48'b100000010010011110000010000110111101100001011010 :
(key == 11'b00001101100) ? 48'b100000010001100011101000000110111010001110000101 :
(key == 11'b00001101101) ? 48'b100000010000101001010100000110110110111011001111 :
(key == 11'b00001101110) ? 48'b100000001111101111000100000110110011101000110100 :
(key == 11'b00001101111) ? 48'b100000001110110100111000000110110000010110111000 :
(key == 11'b00001110000) ? 48'b100000001101111010110100000110101101000101011110 :
(key == 11'b00001110001) ? 48'b100000001101000000110010000110101001110100011011 :
(key == 11'b00001110010) ? 48'b100000001100000110110101000110100110100011110110 :
(key == 11'b00001110011) ? 48'b100000001011001100111110000110100011010011110010 :
(key == 11'b00001110100) ? 48'b100000001010010011001100000110100000000100001010 :
(key == 11'b00001110101) ? 48'b100000001001011001011101000110011100110100111100 :
(key == 11'b00001110110) ? 48'b100000001000011111110100000110011001100110001100 :
(key == 11'b00001110111) ? 48'b100000000111100110010001000110010110010111111101 :
(key == 11'b00001111000) ? 48'b100000000110101100110001000110010011001010000110 :
(key == 11'b00001111001) ? 48'b100000000101110011010111000110001111111100101110 :
(key == 11'b00001111010) ? 48'b100000000100111010000001000110001100101111110010 :
(key == 11'b00001111011) ? 48'b100000000100000000110001000110001001100011010100 :
(key == 11'b00001111100) ? 48'b100000000011000111100110000110000110010111010100 :
(key == 11'b00001111101) ? 48'b100000000010001110011101000110000011001011101010 :
(key == 11'b00001111110) ? 48'b100000000001010101011011000110000000000000100001 :
(key == 11'b00001111111) ? 48'b100000000000011100011110000101111100110101110101 :
(key == 11'b00010000000) ? 48'b011111111111100011100101100101111001101011100110 :
(key == 11'b00010000001) ? 48'b011111111110101010110001000101110110100001101110 :
(key == 11'b00010000010) ? 48'b011111111101110010000001000101110011011000010100 :
(key == 11'b00010000011) ? 48'b011111111100111001010110000101110000001111010110 :
(key == 11'b00010000100) ? 48'b011111111100000000110000100101101101000110110101 :
(key == 11'b00010000101) ? 48'b011111111011001000001111000101101001111110101111 :
(key == 11'b00010000110) ? 48'b011111111010001111110010100101100110110111000101 :
(key == 11'b00010000111) ? 48'b011111111001010111011010000101100011101111110101 :
(key == 11'b00010001000) ? 48'b011111111000011111000111000101100000101001000010 :
(key == 11'b00010001001) ? 48'b011111110111100110111001100101011101100010101110 :
(key == 11'b00010001010) ? 48'b011111110110101110101111000101011010011100101110 :
(key == 11'b00010001011) ? 48'b011111110101110110101001000101010111010111001100 :
(key == 11'b00010001100) ? 48'b011111110100111110101001000101010100010010001000 :
(key == 11'b00010001101) ? 48'b011111110100000110101100000101010001001101011000 :
(key == 11'b00010001110) ? 48'b011111110011001110110100100101001110001001001001 :
(key == 11'b00010001111) ? 48'b011111110010010111000010100101001011000101010111 :
(key == 11'b00010010000) ? 48'b011111110001011111010011100101001000000001111010 :
(key == 11'b00010010001) ? 48'b011111110000100111101010000101000100111110111010 :
(key == 11'b00010010010) ? 48'b011111101111110000000100100101000001111100010101 :
(key == 11'b00010010011) ? 48'b011111101110111000100100100100111110111010001100 :
(key == 11'b00010010100) ? 48'b011111101110000001001000000100111011111000011100 :
(key == 11'b00010010101) ? 48'b011111101101001001110000100100111000110111000101 :
(key == 11'b00010010110) ? 48'b011111101100010010011101000100110101110110001001 :
(key == 11'b00010010111) ? 48'b011111101011011011001111000100110010110101101010 :
(key == 11'b00010011000) ? 48'b011111101010100100000100000100101111110101011111 :
(key == 11'b00010011001) ? 48'b011111101001101100111111000100101100110101110100 :
(key == 11'b00010011010) ? 48'b011111101000110101111110000100101001110110100000 :
(key == 11'b00010011011) ? 48'b011111100111111111000010000100100110110111101001 :
(key == 11'b00010011100) ? 48'b011111100111001000001010100100100011111001001100 :
(key == 11'b00010011101) ? 48'b011111100110010001010111000100100000111011000110 :
(key == 11'b00010011110) ? 48'b011111100101011010100111100100011101111101011011 :
(key == 11'b00010011111) ? 48'b011111100100100011111100000100011011000000000110 :
(key == 11'b00010100000) ? 48'b011111100011101101010110100100011000000011010000 :
(key == 11'b00010100001) ? 48'b011111100010110110110101000100010101000110110010 :
(key == 11'b00010100010) ? 48'b011111100010000000010111000100010010001010101010 :
(key == 11'b00010100011) ? 48'b011111100001001001111110000100001111001111000000 :
(key == 11'b00010100100) ? 48'b011111100000010011101001000100001100010011101011 :
(key == 11'b00010100101) ? 48'b011111011111011101011000100100001001011000110001 :
(key == 11'b00010100110) ? 48'b011111011110100111001100100100000110011110010000 :
(key == 11'b00010100111) ? 48'b011111011101110001000110000100000011100100001011 :
(key == 11'b00010101000) ? 48'b011111011100111011000010000100000000101010011011 :
(key == 11'b00010101001) ? 48'b011111011100000101000011000011111101110001000011 :
(key == 11'b00010101010) ? 48'b011111011011001111001001000011111010111000001000 :
(key == 11'b00010101011) ? 48'b011111011010011001010010100011110111111111100100 :
(key == 11'b00010101100) ? 48'b011111011001100011100001000011110101000111011001 :
(key == 11'b00010101101) ? 48'b011111011000101101110011100011110010001111100111 :
(key == 11'b00010101110) ? 48'b011111010111111000001010000011101111011000001100 :
(key == 11'b00010101111) ? 48'b011111010111000010100101000011101100100001001010 :
(key == 11'b00010110000) ? 48'b011111010110001101000100100011101001101010100000 :
(key == 11'b00010110001) ? 48'b011111010101010111101000100011100110110100010001 :
(key == 11'b00010110010) ? 48'b011111010100100010001111100011100011111110010101 :
(key == 11'b00010110011) ? 48'b011111010011101100111100000011100001001000110100 :
(key == 11'b00010110100) ? 48'b011111010010110111101100100011011110010011101101 :
(key == 11'b00010110101) ? 48'b011111010010000010100001000011011011011110111100 :
(key == 11'b00010110110) ? 48'b011111010001001101011010000011011000101010100100 :
(key == 11'b00010110111) ? 48'b011111010000011000010111100011010101110110100100 :
(key == 11'b00010111000) ? 48'b011111001111100011011001000011010011000010111011 :
(key == 11'b00010111001) ? 48'b011111001110101110011110100011010000001111101011 :
(key == 11'b00010111010) ? 48'b011111001101111001100111000011001101011100101110 :
(key == 11'b00010111011) ? 48'b011111001101000100110101000011001010101010001100 :
(key == 11'b00010111100) ? 48'b011111001100010000001000100011000111111000000110 :
(key == 11'b00010111101) ? 48'b011111001011011011011111000011000101000110010011 :
(key == 11'b00010111110) ? 48'b011111001010100110111001000011000010010100110111 :
(key == 11'b00010111111) ? 48'b011111001001110010010111000010111111100011110010 :
(key == 11'b00011000000) ? 48'b011111001000111101111010000010111100110011000111 :
(key == 11'b00011000001) ? 48'b011111001000001001100001000010111010000010110001 :
(key == 11'b00011000010) ? 48'b011111000111010101001011100010110111010010110001 :
(key == 11'b00011000011) ? 48'b011111000110100000111011000010110100100011001100 :
(key == 11'b00011000100) ? 48'b011111000101101100101110000010110001110011111010 :
(key == 11'b00011000101) ? 48'b011111000100111000100101000010101111000101000000 :
(key == 11'b00011000110) ? 48'b011111000100000100100001000010101100010110011111 :
(key == 11'b00011000111) ? 48'b011111000011010000100000100010101001101000010011 :
(key == 11'b00011001000) ? 48'b011111000010011100100100100010100110111010100000 :
(key == 11'b00011001001) ? 48'b011111000001101000101011100010100100001100111111 :
(key == 11'b00011001010) ? 48'b011111000000110100111000000010100001011111111010 :
(key == 11'b00011001011) ? 48'b011111000000000001000111000010011110110011000111 :
(key == 11'b00011001100) ? 48'b011110111111001101011011100010011100000110101111 :
(key == 11'b00011001101) ? 48'b011110111110011001110011000010011001011010101010 :
(key == 11'b00011001110) ? 48'b011110111101100110001110000010010110101110111010 :
(key == 11'b00011001111) ? 48'b011110111100110010101111000010010100000011100100 :
(key == 11'b00011010000) ? 48'b011110111011111111010011000010010001011000100100 :
(key == 11'b00011010001) ? 48'b011110111011001011111010000010001110101101110111 :
(key == 11'b00011010010) ? 48'b011110111010011000100111000010001100000011100100 :
(key == 11'b00011010011) ? 48'b011110111001100101010110000010001001011001100100 :
(key == 11'b00011010100) ? 48'b011110111000110010001011000010000110101111111110 :
(key == 11'b00011010101) ? 48'b011110110111111111000011000010000100000110101011 :
(key == 11'b00011010110) ? 48'b011110110111001011111110000010000001011101101101 :
(key == 11'b00011010111) ? 48'b011110110110011000111101100001111110110101000100 :
(key == 11'b00011011000) ? 48'b011110110101100110000010000001111100001100110101 :
(key == 11'b00011011001) ? 48'b011110110100110011001001100001111001100100111001 :
(key == 11'b00011011010) ? 48'b011110110100000000010101000001110110111101010010 :
(key == 11'b00011011011) ? 48'b011110110011001101100100000001110100010101111111 :
(key == 11'b00011011100) ? 48'b011110110010011010111000000001110001101111000111 :
(key == 11'b00011011101) ? 48'b011110110001101000001110100001101111001000011111 :
(key == 11'b00011011110) ? 48'b011110110000110101101011000001101100100010010011 :
(key == 11'b00011011111) ? 48'b011110110000000011001010000001101001111100010110 :
(key == 11'b00011100000) ? 48'b011110101111010000101101000001100111010110110010 :
(key == 11'b00011100001) ? 48'b011110101110011110010100000001100100110001100001 :
(key == 11'b00011100010) ? 48'b011110101101101011111110000001100010001100100100 :
(key == 11'b00011100011) ? 48'b011110101100111001101100100001011111100111111101 :
(key == 11'b00011100100) ? 48'b011110101100000111011111100001011101000011101101 :
(key == 11'b00011100101) ? 48'b011110101011010101010110000001011010011111110010 :
(key == 11'b00011100110) ? 48'b011110101010100011010000000001010111111100001010 :
(key == 11'b00011100111) ? 48'b011110101001110001001101100001010101011000110110 :
(key == 11'b00011101000) ? 48'b011110101000111111001111100001010010110101111000 :
(key == 11'b00011101001) ? 48'b011110101000001101010101000001010000010011010000 :
(key == 11'b00011101010) ? 48'b011110100111011011011111000001001101110000111011 :
(key == 11'b00011101011) ? 48'b011110100110101001101011000001001011001110111001 :
(key == 11'b00011101100) ? 48'b011110100101110111111101000001001000101101010001 :
(key == 11'b00011101101) ? 48'b011110100101000110010010000001000110001011111010 :
(key == 11'b00011101110) ? 48'b011110100100010100101010000001000011101010110111 :
(key == 11'b00011101111) ? 48'b011110100011100011000111000001000001001010001011 :
(key == 11'b00011110000) ? 48'b011110100010110001100111000000111110101001110010 :
(key == 11'b00011110001) ? 48'b011110100010000000001011000000111100001001101100 :
(key == 11'b00011110010) ? 48'b011110100001001110110010100000111001101001111010 :
(key == 11'b00011110011) ? 48'b011110100000011101011110100000110111001010011111 :
(key == 11'b00011110100) ? 48'b011110011111101100001101000000110100101011010100 :
(key == 11'b00011110101) ? 48'b011110011110111010111111100000110010001100011111 :
(key == 11'b00011110110) ? 48'b011110011110001001110111000000101111101110000001 :
(key == 11'b00011110111) ? 48'b011110011101011000110000000000101101001111110001 :
(key == 11'b00011111000) ? 48'b011110011100100111101111000000101010110001111011 :
(key == 11'b00011111001) ? 48'b011110011011110110110001000000101000010100010110 :
(key == 11'b00011111010) ? 48'b011110011011000101110101100000100101110111000011 :
(key == 11'b00011111011) ? 48'b011110011010010100111111000000100011011010000110 :
(key == 11'b00011111100) ? 48'b011110011001100100001100000000100000111101011101 :
(key == 11'b00011111101) ? 48'b011110011000110011011100000000011110100001000110 :
(key == 11'b00011111110) ? 48'b011110011000000010101111100000011100000101000010 :
(key == 11'b00011111111) ? 48'b011110010111010010000111000000011001101001010010 :
(key == 11'b00100000000) ? 48'b011110010110100001100010000000010111001101110110 :
(key == 11'b00100000001) ? 48'b011110010101110001000010000000010100110010110001 :
(key == 11'b00100000010) ? 48'b011110010101000000100101000000010010010111111100 :
(key == 11'b00100000011) ? 48'b011110010100010000001011000000001111111101011011 :
(key == 11'b00100000100) ? 48'b011110010011011111110101000000001101100011001100 :
(key == 11'b00100000101) ? 48'b011110010010101111100010000000001011001001010000 :
(key == 11'b00100000110) ? 48'b011110010001111111010011000000001000101111100111 :
(key == 11'b00100000111) ? 48'b011110010001001111001000000000000110010110010011 :
(key == 11'b00100001000) ? 48'b011110010000011111000001000000000011111101010100 :
(key == 11'b00100001001) ? 48'b011110001111101110111100100000000001100100100100 :
(key == 11'b00100001010) ? 48'b011110001110111110111100011111111110011000001111 :
(key == 11'b00100001011) ? 48'b011110001110001110111111011111111001100111111100 :
(key == 11'b00100001100) ? 48'b011110001101011111000101111111110100111000010001 :
(key == 11'b00100001101) ? 48'b011110001100101111001111011111110000001001001000 :
(key == 11'b00100001110) ? 48'b011110001011111111011101111111101011011010101010 :
(key == 11'b00100001111) ? 48'b011110001011001111101111011111100110101100101110 :
(key == 11'b00100010000) ? 48'b011110001010100000000011011111100001111111010011 :
(key == 11'b00100010001) ? 48'b011110001001110000011011011111011101010010100000 :
(key == 11'b00100010010) ? 48'b011110001001000000110111011111011000100110010011 :
(key == 11'b00100010011) ? 48'b011110001000010001010111011111010011111010110010 :
(key == 11'b00100010100) ? 48'b011110000111100001111001011111001111001111101000 :
(key == 11'b00100010101) ? 48'b011110000110110010100000011111001010100101001110 :
(key == 11'b00100010110) ? 48'b011110000110000011001001011111000101111011010000 :
(key == 11'b00100010111) ? 48'b011110000101010011110111011111000001010001111111 :
(key == 11'b00100011000) ? 48'b011110000100100100100111111110111100101001001110 :
(key == 11'b00100011001) ? 48'b011110000011110101011011011110111000000000111111 :
(key == 11'b00100011010) ? 48'b011110000011000110010011111110110011011001011010 :
(key == 11'b00100011011) ? 48'b011110000010010111001111011110101110110010010110 :
(key == 11'b00100011100) ? 48'b011110000001101000001110011110101010001011111001 :
(key == 11'b00100011101) ? 48'b011110000000111001001111011110100101100101111000 :
(key == 11'b00100011110) ? 48'b011110000000001010010101011110100001000000100011 :
(key == 11'b00100011111) ? 48'b011101111111011011011101111110011100011011101101 :
(key == 11'b00100100000) ? 48'b011101111110101100101010011110010111110111011101 :
(key == 11'b00100100001) ? 48'b011101111101111101111010011110010011010011110011 :
(key == 11'b00100100010) ? 48'b011101111101001111001101011110001110110000100101 :
(key == 11'b00100100011) ? 48'b011101111100100000100100011110001010001110000010 :
(key == 11'b00100100100) ? 48'b011101111011110001111110011110000101101100000000 :
(key == 11'b00100100101) ? 48'b011101111011000011011011111110000001001010100010 :
(key == 11'b00100100110) ? 48'b011101111010010100111100011101111100101001100101 :
(key == 11'b00100100111) ? 48'b011101111001100110100000011101111000001001001001 :
(key == 11'b00100101000) ? 48'b011101111000111000001000011101110011101001010111 :
(key == 11'b00100101001) ? 48'b011101111000001001110011011101101111001010000001 :
(key == 11'b00100101010) ? 48'b011101110111011011100010011101101010101011010101 :
(key == 11'b00100101011) ? 48'b011101110110101101010011011101100110001101000101 :
(key == 11'b00100101100) ? 48'b011101110101111111000111011101100001101111010100 :
(key == 11'b00100101101) ? 48'b011101110101010000111111011101011101010010001000 :
(key == 11'b00100101110) ? 48'b011101110100100010111100011101011000110101100111 :
(key == 11'b00100101111) ? 48'b011101110011110100111010111101010100011001100001 :
(key == 11'b00100110000) ? 48'b011101110011000110111101011101001111111110000001 :
(key == 11'b00100110001) ? 48'b011101110010011001000010111101001011100011000000 :
(key == 11'b00100110010) ? 48'b011101110001101011001100011101000111001000100011 :
(key == 11'b00100110011) ? 48'b011101110000111101011001011101000010101110101011 :
(key == 11'b00100110100) ? 48'b011101110000001111101000011100111110010101001110 :
(key == 11'b00100110101) ? 48'b011101101111100001111010011100111001111100010011 :
(key == 11'b00100110110) ? 48'b011101101110110100010001011100110101100011111111 :
(key == 11'b00100110111) ? 48'b011101101110000110101010011100110001001100001000 :
(key == 11'b00100111000) ? 48'b011101101101011001000111111100101100110100111000 :
(key == 11'b00100111001) ? 48'b011101101100101011100111011100101000011110000101 :
(key == 11'b00100111010) ? 48'b011101101011111110001010011100100100000111110000 :
(key == 11'b00100111011) ? 48'b011101101011010000110001011100011111110010000101 :
(key == 11'b00100111100) ? 48'b011101101010100011011011011100011011011100110101 :
(key == 11'b00100111101) ? 48'b011101101001110110000111011100010111001000000100 :
(key == 11'b00100111110) ? 48'b011101101001001000110111111100010010110011111000 :
(key == 11'b00100111111) ? 48'b011101101000011011101011111100001110100000001111 :
(key == 11'b00101000000) ? 48'b011101100111101110100010011100001010001101000010 :
(key == 11'b00101000001) ? 48'b011101100111000001011100011100000101111010010111 :
(key == 11'b00101000010) ? 48'b011101100110010100011001111100000001101000010001 :
(key == 11'b00101000011) ? 48'b011101100101100111011001111011111101010110100111 :
(key == 11'b00101000100) ? 48'b011101100100111010011101011011111001000101011111 :
(key == 11'b00101000101) ? 48'b011101100100001101100100011011110100110100111000 :
(key == 11'b00101000110) ? 48'b011101100011100000101110011011110000100100101110 :
(key == 11'b00101000111) ? 48'b011101100010110011111011011011101100010101001000 :
(key == 11'b00101001000) ? 48'b011101100010000111001011011011101000000101111101 :
(key == 11'b00101001001) ? 48'b011101100001011010011111011011100011110111011010 :
(key == 11'b00101001010) ? 48'b011101100000101101110110011011011111101001010010 :
(key == 11'b00101001011) ? 48'b011101100000000001001111011011011011011011101000 :
(key == 11'b00101001100) ? 48'b011101011111010100101100111011010111001110100011 :
(key == 11'b00101001101) ? 48'b011101011110101000001101011011010011000001111011 :
(key == 11'b00101001110) ? 48'b011101011101111011110000011011001110110101110010 :
(key == 11'b00101001111) ? 48'b011101011101001111010110011011001010101010001000 :
(key == 11'b00101010000) ? 48'b011101011100100011000000011011000110011111000001 :
(key == 11'b00101010001) ? 48'b011101011011110110101101011011000010010100011001 :
(key == 11'b00101010010) ? 48'b011101011011001010011100111010111110001010001011 :
(key == 11'b00101010011) ? 48'b011101011010011110001111111010111010000000100000 :
(key == 11'b00101010100) ? 48'b011101011001110010000101111010110101110111010100 :
(key == 11'b00101010101) ? 48'b011101011001000101111110111010110001101110100101 :
(key == 11'b00101010110) ? 48'b011101011000011001111010111010101101100110010110 :
(key == 11'b00101010111) ? 48'b011101010111101101111011011010101001011110101110 :
(key == 11'b00101011000) ? 48'b011101010111000001111101011010100101010111011010 :
(key == 11'b00101011001) ? 48'b011101010110010110000010011010100001010000100101 :
(key == 11'b00101011010) ? 48'b011101010101101010001011011010011101001010010011 :
(key == 11'b00101011011) ? 48'b011101010100111110010110111010011001000100011111 :
(key == 11'b00101011100) ? 48'b011101010100010010100101011010010100111111001001 :
(key == 11'b00101011101) ? 48'b011101010011100110110111011010010000111010010010 :
(key == 11'b00101011110) ? 48'b011101010010111011001100011010001100110101111000 :
(key == 11'b00101011111) ? 48'b011101010010001111100011111010001000110001111100 :
(key == 11'b00101100000) ? 48'b011101010001100011111111011010000100101110100011 :
(key == 11'b00101100001) ? 48'b011101010000111000011101011010000000101011100011 :
(key == 11'b00101100010) ? 48'b011101010000001100111110011001111100101001000101 :
(key == 11'b00101100011) ? 48'b011101001111100001100011011001111000100111000101 :
(key == 11'b00101100100) ? 48'b011101001110110110001001011001110100100101011010 :
(key == 11'b00101100101) ? 48'b011101001110001010110011011001110000100100010111 :
(key == 11'b00101100110) ? 48'b011101001101011111011111011001101100100011100111 :
(key == 11'b00101100111) ? 48'b011101001100110100010000011001101000100011011111 :
(key == 11'b00101101000) ? 48'b011101001100001001000011011001100100100011110011 :
(key == 11'b00101101001) ? 48'b011101001011011101111001011001100000100100100001 :
(key == 11'b00101101010) ? 48'b011101001010110010110010111001011100100101110001 :
(key == 11'b00101101011) ? 48'b011101001010000111101110011001011000100111011010 :
(key == 11'b00101101100) ? 48'b011101001001011100101101011001010100101001011111 :
(key == 11'b00101101101) ? 48'b011101001000110001101111111001010000101100000111 :
(key == 11'b00101101110) ? 48'b011101001000000110110100011001001100101111001001 :
(key == 11'b00101101111) ? 48'b011101000111011011111100011001001000110010100111 :
(key == 11'b00101110000) ? 48'b011101000110110001000111111001000100110110100111 :
(key == 11'b00101110001) ? 48'b011101000110000110010101011001000000111011000000 :
(key == 11'b00101110010) ? 48'b011101000101011011100110011000111100111111110110 :
(key == 11'b00101110011) ? 48'b011101000100110000111010011000111001000101001001 :
(key == 11'b00101110100) ? 48'b011101000100000110010000011000110101001010110101 :
(key == 11'b00101110101) ? 48'b011101000011011011101001111000110001010001000010 :
(key == 11'b00101110110) ? 48'b011101000010110001000110011000101101010111101100 :
(key == 11'b00101110111) ? 48'b011101000010000110100101011000101001011110101111 :
(key == 11'b00101111000) ? 48'b011101000001011100001000011000100101100110010100 :
(key == 11'b00101111001) ? 48'b011101000000110001101101011000100001101110010000 :
(key == 11'b00101111010) ? 48'b011101000000000111010110011000011101110110101110 :
(key == 11'b00101111011) ? 48'b011100111111011101000000011000011001111111100001 :
(key == 11'b00101111100) ? 48'b011100111110110010101110011000010110001000110100 :
(key == 11'b00101111101) ? 48'b011100111110001000100000011000010010010010101000 :
(key == 11'b00101111110) ? 48'b011100111101011110010011011000001110011100110000 :
(key == 11'b00101111111) ? 48'b011100111100110100001010011000001010100111011001 :
(key == 11'b00110000000) ? 48'b011100111100001010000011011000000110110010011010 :
(key == 11'b00110000001) ? 48'b011100111011011111111111111000000010111101111000 :
(key == 11'b00110000010) ? 48'b011100111010110101111111010111111111001001110010 :
(key == 11'b00110000011) ? 48'b011100111010001100000001010111111011010110001010 :
(key == 11'b00110000100) ? 48'b011100111001100010000101110111110111100010111001 :
(key == 11'b00110000101) ? 48'b011100111000111000001110010111110011110000001001 :
(key == 11'b00110000110) ? 48'b011100111000001110011000010111101111111101110001 :
(key == 11'b00110000111) ? 48'b011100110111100100100110010111101100001011110110 :
(key == 11'b00110001000) ? 48'b011100110110111010110101110111101000011010010010 :
(key == 11'b00110001001) ? 48'b011100110110010001001001010111100100101001001110 :
(key == 11'b00110001010) ? 48'b011100110101100111011111010111100000111000100011 :
(key == 11'b00110001011) ? 48'b011100110100111101110111110111011101001000010100 :
(key == 11'b00110001100) ? 48'b011100110100010100010010110111011001011000011100 :
(key == 11'b00110001101) ? 48'b011100110011101010110001010111010101101001000101 :
(key == 11'b00110001110) ? 48'b011100110011000001010010010111010001111010000110 :
(key == 11'b00110001111) ? 48'b011100110010010111110110010111001110001011100011 :
(key == 11'b00110010000) ? 48'b011100110001101110011101010111001010011101011100 :
(key == 11'b00110010001) ? 48'b011100110001000101000110110111000110101111101100 :
(key == 11'b00110010010) ? 48'b011100110000011011110011010111000011000010011001 :
(key == 11'b00110010011) ? 48'b011100101111110010100011010110111111010101100110 :
(key == 11'b00110010100) ? 48'b011100101111001001010100010110111011101001000101 :
(key == 11'b00110010101) ? 48'b011100101110100000001001010110110111111101000001 :
(key == 11'b00110010110) ? 48'b011100101101110111000000010110110100010001011000 :
(key == 11'b00110010111) ? 48'b011100101101001101111011010110110000100110001010 :
(key == 11'b00110011000) ? 48'b011100101100100100110111110110101100111011010101 :
(key == 11'b00110011001) ? 48'b011100101011111011110110110110101001010000110110 :
(key == 11'b00110011010) ? 48'b011100101011010010111010010110100101100110111100 :
(key == 11'b00110011011) ? 48'b011100101010101001111110010110100001111101010001 :
(key == 11'b00110011100) ? 48'b011100101010000001000110010110011110010100000110 :
(key == 11'b00110011101) ? 48'b011100101001011000010000110110011010101011010001 :
(key == 11'b00110011110) ? 48'b011100101000101111011110110110010111000010111100 :
(key == 11'b00110011111) ? 48'b011100101000000110101110010110010011011010111011 :
(key == 11'b00110100000) ? 48'b011100100111011110000001010110001111110011011001 :
(key == 11'b00110100001) ? 48'b011100100110110101010111010110001100001100001110 :
(key == 11'b00110100010) ? 48'b011100100110001100101110110110001000100101011010 :
(key == 11'b00110100011) ? 48'b011100100101100100001010010110000100111111000110 :
(key == 11'b00110100100) ? 48'b011100100100111011101000010110000001011001001000 :
(key == 11'b00110100101) ? 48'b011100100100010011001000010101111101110011100001 :
(key == 11'b00110100110) ? 48'b011100100011101010101011010101111010001110010110 :
(key == 11'b00110100111) ? 48'b011100100011000010010001010101110110101001100101 :
(key == 11'b00110101000) ? 48'b011100100010011001111001010101110011000101001100 :
(key == 11'b00110101001) ? 48'b011100100001110001100100010101101111100001001110 :
(key == 11'b00110101010) ? 48'b011100100001001001010010010101101011111101100110 :
(key == 11'b00110101011) ? 48'b011100100000100001000001110101101000011010010101 :
(key == 11'b00110101100) ? 48'b011100011111111000110110010101100100110111101000 :
(key == 11'b00110101101) ? 48'b011100011111010000101011010101100001010101001000 :
(key == 11'b00110101110) ? 48'b011100011110101000100011010101011101110011000100 :
(key == 11'b00110101111) ? 48'b011100011110000000011110010101011010010001011010 :
(key == 11'b00110110000) ? 48'b011100011101011000011011010101010110110000000111 :
(key == 11'b00110110001) ? 48'b011100011100110000011100010101010011001111010011 :
(key == 11'b00110110010) ? 48'b011100011100001000011110110101001111101110110001 :
(key == 11'b00110110011) ? 48'b011100011011100000100101010101001100001110101111 :
(key == 11'b00110110100) ? 48'b011100011010111000101100110101001000101110111110 :
(key == 11'b00110110101) ? 48'b011100011010010000110111010101000101001111101000 :
(key == 11'b00110110110) ? 48'b011100011001101001000100010101000001110000101000 :
(key == 11'b00110110111) ? 48'b011100011001000001010100010100111110010010000100 :
(key == 11'b00110111000) ? 48'b011100011000011001100111010100111010110011111001 :
(key == 11'b00110111001) ? 48'b011100010111110001111100110100110111010110000101 :
(key == 11'b00110111010) ? 48'b011100010111001010010100010100110011111000100111 :
(key == 11'b00110111011) ? 48'b011100010110100010101110110100110000011011100011 :
(key == 11'b00110111100) ? 48'b011100010101111011001011010100101100111110110110 :
(key == 11'b00110111101) ? 48'b011100010101010011101011010100101001100010100011 :
(key == 11'b00110111110) ? 48'b011100010100101100001101010100100110000110100110 :
(key == 11'b00110111111) ? 48'b011100010100000100110010010100100010101011000100 :
(key == 11'b00111000000) ? 48'b011100010011011101011001010100011111001111110111 :
(key == 11'b00111000001) ? 48'b011100010010110110000011010100011011110101000000 :
(key == 11'b00111000010) ? 48'b011100010010001110101111010100011000011010100100 :
(key == 11'b00111000011) ? 48'b011100010001100111011111010100010101000000100010 :
(key == 11'b00111000100) ? 48'b011100010001000000010000010100010001100110110010 :
(key == 11'b00111000101) ? 48'b011100010000011001000011010100001110001101010111 :
(key == 11'b00111000110) ? 48'b011100001111110001111010010100001010110100011010 :
(key == 11'b00111000111) ? 48'b011100001111001010110100010100000111011011111000 :
(key == 11'b00111001000) ? 48'b011100001110100011101111010100000100000011100100 :
(key == 11'b00111001001) ? 48'b011100001101111100101101010100000000101011101101 :
(key == 11'b00111001010) ? 48'b011100001101010101101111010011111101010100010000 :
(key == 11'b00111001011) ? 48'b011100001100101110110010010011111001111101000101 :
(key == 11'b00111001100) ? 48'b011100001100000111111000010011110110100110010100 :
(key == 11'b00111001101) ? 48'b011100001011100000111111010011110011001111110100 :
(key == 11'b00111001110) ? 48'b011100001010111010001010010011101111111001101110 :
(key == 11'b00111001111) ? 48'b011100001010010011011000010011101100100100000110 :
(key == 11'b00111010000) ? 48'b011100001001101100101000010011101001001110101111 :
(key == 11'b00111010001) ? 48'b011100001001000101111010010011100101111001101110 :
(key == 11'b00111010010) ? 48'b011100001000011111001111010011100010100101000110 :
(key == 11'b00111010011) ? 48'b011100000111111000100111010011011111010000111000 :
(key == 11'b00111010100) ? 48'b011100000111010001111111110011011011111100111000 :
(key == 11'b00111010101) ? 48'b011100000110101011011100010011011000101001010101 :
(key == 11'b00111010110) ? 48'b011100000110000100111011110011010101010110001011 :
(key == 11'b00111010111) ? 48'b011100000101011110011100110011010010000011010011 :
(key == 11'b00111011000) ? 48'b011100000100111000000000010011001110110000110000 :
(key == 11'b00111011001) ? 48'b011100000100010001100110010011001011011110100111 :
(key == 11'b00111011010) ? 48'b011100000011101011001110110011001000001100110010 :
(key == 11'b00111011011) ? 48'b011100000011000100111010010011000100111011011000 :
(key == 11'b00111011100) ? 48'b011100000010011110100111010011000001101010001110 :
(key == 11'b00111011101) ? 48'b011100000001111000010111010010111110011001011110 :
(key == 11'b00111011110) ? 48'b011100000001010010001001010010111011001001000010 :
(key == 11'b00111011111) ? 48'b011100000000101011111110110010110111111001000000 :
(key == 11'b00111100000) ? 48'b011100000000000101110101010010110100101001001111 :
(key == 11'b00111100001) ? 48'b011011111111011111110000010010110001011001111100 :
(key == 11'b00111100010) ? 48'b011011111110111001101011010010101110001010110100 :
(key == 11'b00111100011) ? 48'b011011111110010011101010010010101010111100001011 :
(key == 11'b00111100100) ? 48'b011011111101101101101011010010100111101101110110 :
(key == 11'b00111100101) ? 48'b011011111101000111101111010010100100011111110110 :
(key == 11'b00111100110) ? 48'b011011111100100001110100110010100001010010001100 :
(key == 11'b00111100111) ? 48'b011011111011111011111100110010011110000100110110 :
(key == 11'b00111101000) ? 48'b011011111011010110000111110010011010110111111001 :
(key == 11'b00111101001) ? 48'b011011111010110000010101010010010111101011010000 :
(key == 11'b00111101010) ? 48'b011011111010001010100011110010010100011110111001 :
(key == 11'b00111101011) ? 48'b011011111001100100110110010010010001010010111111 :
(key == 11'b00111101100) ? 48'b011011111000111111001010010010001110000111010101 :
(key == 11'b00111101101) ? 48'b011011111000011001100000010010001010111100000000 :
(key == 11'b00111101110) ? 48'b011011110111110011111001110010000111110001000100 :
(key == 11'b00111101111) ? 48'b011011110111001110010101010010000100100110011100 :
(key == 11'b00111110000) ? 48'b011011110110101000110010010010000001011100000101 :
(key == 11'b00111110001) ? 48'b011011110110000011010011010001111110010010001011 :
(key == 11'b00111110010) ? 48'b011011110101011101110110010001111011001000100101 :
(key == 11'b00111110011) ? 48'b011011110100111000011010010001110111111111010000 :
(key == 11'b00111110100) ? 48'b011011110100010011000010010001110100110110010100 :
(key == 11'b00111110101) ? 48'b011011110011101101101011010001110001101101101000 :
(key == 11'b00111110110) ? 48'b011011110011001000010111010001101110100101010100 :
(key == 11'b00111110111) ? 48'b011011110010100011000100010001101011011101010010 :
(key == 11'b00111111000) ? 48'b011011110001111101110101010001101000010101100111 :
(key == 11'b00111111001) ? 48'b011011110001011000101000010001100101001110010101 :
(key == 11'b00111111010) ? 48'b011011110000110011011110010001100010000111010111 :
(key == 11'b00111111011) ? 48'b011011110000001110010101010001011111000000101010 :
(key == 11'b00111111100) ? 48'b011011101111101001001111110001011011111010010101 :
(key == 11'b00111111101) ? 48'b011011101111000100001011010001011000110100010000 :
(key == 11'b00111111110) ? 48'b011011101110011111001001010001010101101110100000 :
(key == 11'b00111111111) ? 48'b011011101101111010001011010001010010101001001011 :
(key == 11'b01000000000) ? 48'b011011101101010101001110010001001111100100000111 :
(key == 11'b01000000001) ? 48'b011011101100110000010011010001001100011111010011 :
(key == 11'b01000000010) ? 48'b011011101100001011011011110001001001011010111100 :
(key == 11'b01000000011) ? 48'b011011101011100110100101110001000110010110110100 :
(key == 11'b01000000100) ? 48'b011011101011000001110010010001000011010011000001 :
(key == 11'b01000000101) ? 48'b011011101010011101000000010001000000001111100010 :
(key == 11'b01000000110) ? 48'b011011101001111000010001010000111101001100010110 :
(key == 11'b01000000111) ? 48'b011011101001010011100100010000111010001001011111 :
(key == 11'b01000001000) ? 48'b011011101000101110111010010000110111000111000000 :
(key == 11'b01000001001) ? 48'b011011101000001010010010010000110100000100110101 :
(key == 11'b01000001010) ? 48'b011011100111100101101100010000110001000010111010 :
(key == 11'b01000001011) ? 48'b011011100111000001001000010000101110000001010010 :
(key == 11'b01000001100) ? 48'b011011100110011100100111010000101011000000000011 :
(key == 11'b01000001101) ? 48'b011011100101111000000111110000100111111111000100 :
(key == 11'b01000001110) ? 48'b011011100101010011101011010000100100111110011100 :
(key == 11'b01000001111) ? 48'b011011100100101111010001010000100001111110001000 :
(key == 11'b01000010000) ? 48'b011011100100001010111000010000011110111110000100 :
(key == 11'b01000010001) ? 48'b011011100011100110100010010000011011111110011000 :
(key == 11'b01000010010) ? 48'b011011100011000010001110010000011000111110111100 :
(key == 11'b01000010011) ? 48'b011011100010011101111101010000010101111111110111 :
(key == 11'b01000010100) ? 48'b011011100001111001101101010000010011000001000010 :
(key == 11'b01000010101) ? 48'b011011100001010101100000010000010000000010100100 :
(key == 11'b01000010110) ? 48'b011011100000110001010101010000001101000100010111 :
(key == 11'b01000010111) ? 48'b011011100000001101001101010000001010000110100001 :
(key == 11'b01000011000) ? 48'b011011011111101001000110010000000111001000111010 :
(key == 11'b01000011001) ? 48'b011011011111000101000001110000000100001011101000 :
(key == 11'b01000011010) ? 48'b011011011110100001000000010000000001001110101100 :
(key == 11'b01000011011) ? 48'b011011011101111101000000001111111110010010000000 :
(key == 11'b01000011100) ? 48'b011011011101011001000010001111111011010101101000 :
(key == 11'b01000011101) ? 48'b011011011100110101000110001111111000011001100000 :
(key == 11'b01000011110) ? 48'b011011011100010001001101101111110101011101110010 :
(key == 11'b01000011111) ? 48'b011011011011101101010110101111110010100010010101 :
(key == 11'b01000100000) ? 48'b011011011011001001100010001111101111100111001010 :
(key == 11'b01000100001) ? 48'b011011011010100101101111001111101100101100010011 :
(key == 11'b01000100010) ? 48'b011011011010000001111111001111101001110001101111 :
(key == 11'b01000100011) ? 48'b011011011001011110010000001111100110110111011011 :
(key == 11'b01000100100) ? 48'b011011011000111010100100101111100011111101011110 :
(key == 11'b01000100101) ? 48'b011011011000010110111010001111100001000011110000 :
(key == 11'b01000100110) ? 48'b011011010111110011010011001111011110001010011010 :
(key == 11'b01000100111) ? 48'b011011010111001111101101001111011011010001010010 :
(key == 11'b01000101000) ? 48'b011011010110101100001010001111011000011000011110 :
(key == 11'b01000101001) ? 48'b011011010110001000101000101111010101011111111101 :
(key == 11'b01000101010) ? 48'b011011010101100101001001101111010010100111110000 :
(key == 11'b01000101011) ? 48'b011011010101000001101101001111001111101111110110 :
(key == 11'b01000101100) ? 48'b011011010100011110010001101111001100111000001010 :
(key == 11'b01000101101) ? 48'b011011010011111010111001001111001010000000110110 :
(key == 11'b01000101110) ? 48'b011011010011010111100010101111000111001001110001 :
(key == 11'b01000101111) ? 48'b011011010010110100001111001111000100010011000010 :
(key == 11'b01000110000) ? 48'b011011010010010000111101001111000001011100101000 :
(key == 11'b01000110001) ? 48'b011011010001101101101101001110111110100110011100 :
(key == 11'b01000110010) ? 48'b011011010001001010011111001110111011110000011111 :
(key == 11'b01000110011) ? 48'b011011010000100111010011001110111000111010111000 :
(key == 11'b01000110100) ? 48'b011011010000000100001001001110110110000101100010 :
(key == 11'b01000110101) ? 48'b011011001111100001000001101110110011010000011101 :
(key == 11'b01000110110) ? 48'b011011001110111101111101001110110000011011110000 :
(key == 11'b01000110111) ? 48'b011011001110011010111001101110101101100111010010 :
(key == 11'b01000111000) ? 48'b011011001101110111111000101110101010110011000110 :
(key == 11'b01000111001) ? 48'b011011001101010100111001001110100111111111001001 :
(key == 11'b01000111010) ? 48'b011011001100110001111100101110100101001011100011 :
(key == 11'b01000111011) ? 48'b011011001100001111000001101110100010011000001100 :
(key == 11'b01000111100) ? 48'b011011001011101100001000001110011111100101000100 :
(key == 11'b01000111101) ? 48'b011011001011001001010010001110011100110010010110 :
(key == 11'b01000111110) ? 48'b011011001010100110011110001110011001111111110111 :
(key == 11'b01000111111) ? 48'b011011001010000011101010101110010111001101100100 :
(key == 11'b01001000000) ? 48'b011011001001100000111011001110010100011011101010 :
(key == 11'b01001000001) ? 48'b011011001000111110001100001110010001101001111011 :
(key == 11'b01001000010) ? 48'b011011001000011011100000001110001110111000100011 :
(key == 11'b01001000011) ? 48'b011011000111111000110110001110001100000111011101 :
(key == 11'b01001000100) ? 48'b011011000111010110001110001110001001010110100110 :
(key == 11'b01001000101) ? 48'b011011000110110011101000001110000110100110000010 :
(key == 11'b01001000110) ? 48'b011011000110010001000100001110000011110101110000 :
(key == 11'b01001000111) ? 48'b011011000101101110100010001110000001000101101100 :
(key == 11'b01001001000) ? 48'b011011000101001100000010001101111110010101111100 :
(key == 11'b01001001001) ? 48'b011011000100101001100101001101111011100110100010 :
(key == 11'b01001001010) ? 48'b011011000100000111001000101101111000110111010010 :
(key == 11'b01001001011) ? 48'b011011000011100100101111001101110110001000011001 :
(key == 11'b01001001100) ? 48'b011011000011000010010111101101110011011001101110 :
(key == 11'b01001001101) ? 48'b011011000010100000000010001101110000101011010101 :
(key == 11'b01001001110) ? 48'b011011000001111101101111001101101101111101001111 :
(key == 11'b01001001111) ? 48'b011011000001011011011110001101101011001111011011 :
(key == 11'b01001010000) ? 48'b011011000000111001001101101101101000100001110010 :
(key == 11'b01001010001) ? 48'b011011000000010111000000001101100101110100011110 :
(key == 11'b01001010010) ? 48'b011010111111110100110101001101100011000111011110 :
(key == 11'b01001010011) ? 48'b011010111111010010101100001101100000011010101100 :
(key == 11'b01001010100) ? 48'b011010111110110000100100101101011101101110001011 :
(key == 11'b01001010101) ? 48'b011010111110001110011111101101011011000001111110 :
(key == 11'b01001010110) ? 48'b011010111101101100011100001101011000010101111110 :
(key == 11'b01001010111) ? 48'b011010111101001010011011001101010101101010010000 :
(key == 11'b01001011000) ? 48'b011010111100101000011100001101010010111110110100 :
(key == 11'b01001011001) ? 48'b011010111100000110011110001101010000010011100111 :
(key == 11'b01001011010) ? 48'b011010111011100100100011001101001101101000101100 :
(key == 11'b01001011011) ? 48'b011010111011000010101010001101001010111110000011 :
(key == 11'b01001011100) ? 48'b011010111010100000110010101101001000010011101001 :
(key == 11'b01001011101) ? 48'b011010111001111110111101001101000101101001100000 :
(key == 11'b01001011110) ? 48'b011010111001011101001010001101000010111111101001 :
(key == 11'b01001011111) ? 48'b011010111000111011011001001101000000010110000001 :
(key == 11'b01001100000) ? 48'b011010111000011001101001101100111101101100101010 :
(key == 11'b01001100001) ? 48'b011010110111110111111100001100111011000011100010 :
(key == 11'b01001100010) ? 48'b011010110111010110010000001100111000011010101011 :
(key == 11'b01001100011) ? 48'b011010110110110100100111001100110101110010000110 :
(key == 11'b01001100100) ? 48'b011010110110010011000000001100110011001001110100 :
(key == 11'b01001100101) ? 48'b011010110101110001011010101100110000100001101111 :
(key == 11'b01001100110) ? 48'b011010110101001111110111001100101101111001111100 :
(key == 11'b01001100111) ? 48'b011010110100101110010110001100101011010010011011 :
(key == 11'b01001101000) ? 48'b011010110100001100110110001100101000101011000100 :
(key == 11'b01001101001) ? 48'b011010110011101011011001001100100110000100000011 :
(key == 11'b01001101010) ? 48'b011010110011001001111110001100100011011101010011 :
(key == 11'b01001101011) ? 48'b011010110010101000100100001100100000110110110010 :
(key == 11'b01001101100) ? 48'b011010110010000111001100001100011110010000011110 :
(key == 11'b01001101101) ? 48'b011010110001100101110110001100011011101010011000 :
(key == 11'b01001101110) ? 48'b011010110001000100100010001100011001000100101000 :
(key == 11'b01001101111) ? 48'b011010110000100011010001001100010110011111001010 :
(key == 11'b01001110000) ? 48'b011010110000000010000001001100010011111001111001 :
(key == 11'b01001110001) ? 48'b011010101111100000110011001100010001010100110110 :
(key == 11'b01001110010) ? 48'b011010101110111111100110001100001110110000000000 :
(key == 11'b01001110011) ? 48'b011010101110011110011101001100001100001011100101 :
(key == 11'b01001110100) ? 48'b011010101101111101010101001100001001100111010010 :
(key == 11'b01001110101) ? 48'b011010101101011100001110001100000111000011001111 :
(key == 11'b01001110110) ? 48'b011010101100111011001010001100000100011111011100 :
(key == 11'b01001110111) ? 48'b011010101100011010000111101100000001111011111010 :
(key == 11'b01001111000) ? 48'b011010101011111001000111001011111111011000100111 :
(key == 11'b01001111001) ? 48'b011010101011011000001000001011111100110101100101 :
(key == 11'b01001111010) ? 48'b011010101010110111001100001011111010010010110100 :
(key == 11'b01001111011) ? 48'b011010101010010110010001001011110111110000010010 :
(key == 11'b01001111100) ? 48'b011010101001110101011000001011110101001101111100 :
(key == 11'b01001111101) ? 48'b011010101001010100100001001011110010101011111000 :
(key == 11'b01001111110) ? 48'b011010101000110011101100001011110000001010000110 :
(key == 11'b01001111111) ? 48'b011010101000010010111010001011101101101000100100 :
(key == 11'b01010000000) ? 48'b011010100111110010000111001011101011000111001001 :
(key == 11'b01010000001) ? 48'b011010100111010001011000101011101000100110000111 :
(key == 11'b01010000010) ? 48'b011010100110110000101010101011100110000101001110 :
(key == 11'b01010000011) ? 48'b011010100110001111111111101011100011100100101011 :
(key == 11'b01010000100) ? 48'b011010100101101111010110001011100001000100010101 :
(key == 11'b01010000101) ? 48'b011010100101001110101101001011011110100100001000 :
(key == 11'b01010000110) ? 48'b011010100100101110000111101011011100000100010001 :
(key == 11'b01010000111) ? 48'b011010100100001101100100001011011001100100101011 :
(key == 11'b01010001000) ? 48'b011010100011101101000010001011010111000101010010 :
(key == 11'b01010001001) ? 48'b011010100011001100100001001011010100100110000011 :
(key == 11'b01010001010) ? 48'b011010100010101100000010001011010010000111000101 :
(key == 11'b01010001011) ? 48'b011010100010001011100110001011001111101000011100 :
(key == 11'b01010001100) ? 48'b011010100001101011001011001011001101001010000000 :
(key == 11'b01010001101) ? 48'b011010100001001010110010001011001010101011110010 :
(key == 11'b01010001110) ? 48'b011010100000101010011011101011001000001101110100 :
(key == 11'b01010001111) ? 48'b011010100000001010000110001011000101110000000100 :
(key == 11'b01010010000) ? 48'b011010011111101001110010001011000011010010011110 :
(key == 11'b01010010001) ? 48'b011010011111001001100001001011000000110101010000 :
(key == 11'b01010010010) ? 48'b011010011110101001010001001010111110011000001011 :
(key == 11'b01010010011) ? 48'b011010011110001001000011001010111011111011011000 :
(key == 11'b01010010100) ? 48'b011010011101101000110111001010111001011110110001 :
(key == 11'b01010010101) ? 48'b011010011101001000101101001010110111000010011100 :
(key == 11'b01010010110) ? 48'b011010011100101000100100101010110100100110010100 :
(key == 11'b01010010111) ? 48'b011010011100001000011110001010110010001010011100 :
(key == 11'b01010011000) ? 48'b011010011011101000011001001010101111101110101110 :
(key == 11'b01010011001) ? 48'b011010011011001000010110001010101101010011010101 :
(key == 11'b01010011010) ? 48'b011010011010101000010110001010101010111000001100 :
(key == 11'b01010011011) ? 48'b011010011010001000010110101010101000011101001110 :
(key == 11'b01010011100) ? 48'b011010011001101000011001001010100110000010011111 :
(key == 11'b01010011101) ? 48'b011010011001001000011101101010100011100111111110 :
(key == 11'b01010011110) ? 48'b011010011000101000100011001010100001001101101010 :
(key == 11'b01010011111) ? 48'b011010011000001000101011001010011110110011100110 :
(key == 11'b01010100000) ? 48'b011010010111101000110101001010011100011001110000 :
(key == 11'b01010100001) ? 48'b011010010111001001000001001010011010000000001110 :
(key == 11'b01010100010) ? 48'b011010010110101001001110001010010111100110110010 :
(key == 11'b01010100011) ? 48'b011010010110001001011101001010010101001101101010 :
(key == 11'b01010100100) ? 48'b011010010101101001101110001010010010110100101111 :
(key == 11'b01010100101) ? 48'b011010010101001010000001001010010000011100000001 :
(key == 11'b01010100110) ? 48'b011010010100101010010101101010001110000011100011 :
(key == 11'b01010100111) ? 48'b011010010100001010101100101010001011101011010110 :
(key == 11'b01010101000) ? 48'b011010010011101011000100001010001001010011010010 :
(key == 11'b01010101001) ? 48'b011010010011001011011101101010000110111011011100 :
(key == 11'b01010101010) ? 48'b011010010010101011111010001010000100100011111010 :
(key == 11'b01010101011) ? 48'b011010010010001100010111001010000010001100100000 :
(key == 11'b01010101100) ? 48'b011010010001101100110111001001111111110101011011 :
(key == 11'b01010101101) ? 48'b011010010001001101010111101001111101011110011110 :
(key == 11'b01010101110) ? 48'b011010010000101101111010101001111011000111110011 :
(key == 11'b01010101111) ? 48'b011010010000001110011111001001111000110001010101 :
(key == 11'b01010110000) ? 48'b011010001111101111000101001001110110011011000010 :
(key == 11'b01010110001) ? 48'b011010001111001111101100101001110100000100111101 :
(key == 11'b01010110010) ? 48'b011010001110110000010110001001110001101111001000 :
(key == 11'b01010110011) ? 48'b011010001110010001000010001001101111011001100100 :
(key == 11'b01010110100) ? 48'b011010001101110001110000001001101101000100001100 :
(key == 11'b01010110101) ? 48'b011010001101010010011111001001101010101111000010 :
(key == 11'b01010110110) ? 48'b011010001100110011010000001001101000011010000110 :
(key == 11'b01010110111) ? 48'b011010001100010100000011001001100110000101011000 :
(key == 11'b01010111000) ? 48'b011010001011110100110111001001100011110000111000 :
(key == 11'b01010111001) ? 48'b011010001011010101101101001001100001011100100011 :
(key == 11'b01010111010) ? 48'b011010001010110110100100001001011111001000011011 :
(key == 11'b01010111011) ? 48'b011010001010010111011101101001011100110100100011 :
(key == 11'b01010111100) ? 48'b011010001001111000011001001001011010100000111011 :
(key == 11'b01010111101) ? 48'b011010001001011001010110001001011000001101011100 :
(key == 11'b01010111110) ? 48'b011010001000111010010100101001010101111010001110 :
(key == 11'b01010111111) ? 48'b011010001000011011010101001001010011100111001100 :
(key == 11'b01011000000) ? 48'b011010000111111100011000001001010001010100011110 :
(key == 11'b01011000001) ? 48'b011010000111011101011011001001001111000001110101 :
(key == 11'b01011000010) ? 48'b011010000110111110100000001001001100101111011001 :
(key == 11'b01011000011) ? 48'b011010000110011111101000001001001010011101010000 :
(key == 11'b01011000100) ? 48'b011010000110000000110001001001001000001011010100 :
(key == 11'b01011000101) ? 48'b011010000101100001111100001001000101111001100100 :
(key == 11'b01011000110) ? 48'b011010000101000011001000001001000011101000000001 :
(key == 11'b01011000111) ? 48'b011010000100100100010110001001000001010110101010 :
(key == 11'b01011001000) ? 48'b011010000100000101100110001000111111000101100100 :
(key == 11'b01011001001) ? 48'b011010000011100110110111001000111100110100101001 :
(key == 11'b01011001010) ? 48'b011010000011001000001011001000111010100011111111 :
(key == 11'b01011001011) ? 48'b011010000010101001011111101000111000010011011101 :
(key == 11'b01011001100) ? 48'b011010000010001010110110001000110110000011001100 :
(key == 11'b01011001101) ? 48'b011010000001101100001110101000110011110011000110 :
(key == 11'b01011001110) ? 48'b011010000001001101101001001000110001100011010001 :
(key == 11'b01011001111) ? 48'b011010000000101111000100001000101111010011100100 :
(key == 11'b01011010000) ? 48'b011010000000010000100010001000101101000100001000 :
(key == 11'b01011010001) ? 48'b011001111111110010000001001000101010110100110111 :
(key == 11'b01011010010) ? 48'b011001111111010011100001001000101000100101110011 :
(key == 11'b01011010011) ? 48'b011001111110110101000100001000100110010110111110 :
(key == 11'b01011010100) ? 48'b011001111110010110100111101000100100001000010011 :
(key == 11'b01011010101) ? 48'b011001111101111000001110001000100001111001111010 :
(key == 11'b01011010110) ? 48'b011001111101011001110101001000011111101011101011 :
(key == 11'b01011010111) ? 48'b011001111100111011011110001000011101011101100111 :
(key == 11'b01011011000) ? 48'b011001111100011101001001001000011011001111110100 :
(key == 11'b01011011001) ? 48'b011001111011111110110101101000011001000010001100 :
(key == 11'b01011011010) ? 48'b011001111011100000100100001000010110110100110100 :
(key == 11'b01011011011) ? 48'b011001111011000010010011001000010100100111100010 :
(key == 11'b01011011100) ? 48'b011001111010100100000101001000010010011010100010 :
(key == 11'b01011011101) ? 48'b011001111010000101111000001000010000001101101110 :
(key == 11'b01011011110) ? 48'b011001111001100111101101001000001110000001000111 :
(key == 11'b01011011111) ? 48'b011001111001001001100010001000001011110100101000 :
(key == 11'b01011100000) ? 48'b011001111000101011011011001000001001101000011101 :
(key == 11'b01011100001) ? 48'b011001111000001101010100001000000111011100011010 :
(key == 11'b01011100010) ? 48'b011001110111101111001111101000000101010000100110 :
(key == 11'b01011100011) ? 48'b011001110111010001001100101000000011000100111111 :
(key == 11'b01011100100) ? 48'b011001110110110011001011001000000000111001100100 :
(key == 11'b01011100101) ? 48'b011001110110010101001011000111111110101110010100 :
(key == 11'b01011100110) ? 48'b011001110101110111001100100111111100100011010001 :
(key == 11'b01011100111) ? 48'b011001110101011001010000000111111010011000011101 :
(key == 11'b01011101000) ? 48'b011001110100111011010101100111111000001101110101 :
(key == 11'b01011101001) ? 48'b011001110100011101011011100111110110000011010101 :
(key == 11'b01011101010) ? 48'b011001110011111111100100000111110011111001000101 :
(key == 11'b01011101011) ? 48'b011001110011100001101101100111110001101111000001 :
(key == 11'b01011101100) ? 48'b011001110011000011111001000111101111100101001001 :
(key == 11'b01011101101) ? 48'b011001110010100110000110000111101101011011100000 :
(key == 11'b01011101110) ? 48'b011001110010001000010101000111101011010010000011 :
(key == 11'b01011101111) ? 48'b011001110001101010100110000111101001001000110010 :
(key == 11'b01011110000) ? 48'b011001110001001100110111000111100110111111101001 :
(key == 11'b01011110001) ? 48'b011001110000101111001011000111100100110110110100 :
(key == 11'b01011110010) ? 48'b011001110000010001100000000111100010101110000110 :
(key == 11'b01011110011) ? 48'b011001101111110011110111100111100000100101101000 :
(key == 11'b01011110100) ? 48'b011001101111010110001111100111011110011101010010 :
(key == 11'b01011110101) ? 48'b011001101110111000101001000111011100010101001000 :
(key == 11'b01011110110) ? 48'b011001101110011011000101000111011010001101001101 :
(key == 11'b01011110111) ? 48'b011001101101111101100011000111011000000101100001 :
(key == 11'b01011111000) ? 48'b011001101101100000000001000111010101111101111011 :
(key == 11'b01011111001) ? 48'b011001101101000010100001000111010011110110100011 :
(key == 11'b01011111010) ? 48'b011001101100100101000011000111010001101111010111 :
(key == 11'b01011111011) ? 48'b011001101100000111100111000111001111101000011010 :
(key == 11'b01011111100) ? 48'b011001101011101010001011100111001101100001100110 :
(key == 11'b01011111101) ? 48'b011001101011001100110010000111001011011010111101 :
(key == 11'b01011111110) ? 48'b011001101010101111011010000111001001010100100100 :
(key == 11'b01011111111) ? 48'b011001101010010010000100000111000111001110010110 :
(key == 11'b01100000000) ? 48'b011001101001110100110000000111000101001000010100 :
(key == 11'b01100000001) ? 48'b011001101001010111011101000111000011000010011101 :
(key == 11'b01100000010) ? 48'b011001101000111010001010100111000000111100101110 :
(key == 11'b01100000011) ? 48'b011001101000011100111010100110111110110111001111 :
(key == 11'b01100000100) ? 48'b011001100111111111101101000110111100110001111111 :
(key == 11'b01100000101) ? 48'b011001100111100010100000000110111010101100110110 :
(key == 11'b01100000110) ? 48'b011001100111000101010101000110111000100111111101 :
(key == 11'b01100000111) ? 48'b011001100110101000001011000110110110100011001100 :
(key == 11'b01100001000) ? 48'b011001100110001011000010100110110100011110100111 :
(key == 11'b01100001001) ? 48'b011001100101101101111100000110110010011010010000 :
(key == 11'b01100001010) ? 48'b011001100101010000110111100110110000010110000101 :
(key == 11'b01100001011) ? 48'b011001100100110011110011100110101110010010000010 :
(key == 11'b01100001100) ? 48'b011001100100010110110010000110101100001110001110 :
(key == 11'b01100001101) ? 48'b011001100011111001110001000110101010001010100010 :
(key == 11'b01100001110) ? 48'b011001100011011100110011000110101000000111001000 :
(key == 11'b01100001111) ? 48'b011001100010111111110101000110100110000011110011 :
(key == 11'b01100010000) ? 48'b011001100010100010111001000110100100000000101101 :
(key == 11'b01100010001) ? 48'b011001100010000101111111100110100001111101110101 :
(key == 11'b01100010010) ? 48'b011001100001101001000111000110011111111011000110 :
(key == 11'b01100010011) ? 48'b011001100001001100001111000110011101111000011111 :
(key == 11'b01100010100) ? 48'b011001100000101111011010000110011011110110001010 :
(key == 11'b01100010101) ? 48'b011001100000010010100101100110011001110011111100 :
(key == 11'b01100010110) ? 48'b011001011111110101110011000110010111110001111010 :
(key == 11'b01100010111) ? 48'b011001011111011001000001100110010101110000000100 :
(key == 11'b01100011000) ? 48'b011001011110111100010010000110010011101110011001 :
(key == 11'b01100011001) ? 48'b011001011110011111100100000110010001101100111100 :
(key == 11'b01100011010) ? 48'b011001011110000010111000000110001111101011101011 :
(key == 11'b01100011011) ? 48'b011001011101100110001101000110001101101010100010 :
(key == 11'b01100011100) ? 48'b011001011101001001100011000110001011101001100100 :
(key == 11'b01100011101) ? 48'b011001011100101100111011000110001001101000110010 :
(key == 11'b01100011110) ? 48'b011001011100010000010101000110000111101000001110 :
(key == 11'b01100011111) ? 48'b011001011011110011110000000110000101100111110010 :
(key == 11'b01100100000) ? 48'b011001011011010111001101000110000011100111100100 :
(key == 11'b01100100001) ? 48'b011001011010111010101010000110000001100111011011 :
(key == 11'b01100100010) ? 48'b011001011010011110001010000101111111100111100100 :
(key == 11'b01100100011) ? 48'b011001011010000001101011000101111101100111111000 :
(key == 11'b01100100100) ? 48'b011001011001100101001101100101111011101000010100 :
(key == 11'b01100100101) ? 48'b011001011001001000110001000101111001101000111100 :
(key == 11'b01100100110) ? 48'b011001011000101100010111000101110111101001110001 :
(key == 11'b01100100111) ? 48'b011001011000001111111110000101110101101010101111 :
(key == 11'b01100101000) ? 48'b011001010111110011100110000101110011101011110111 :
(key == 11'b01100101001) ? 48'b011001010111010111010001000101110001101101001110 :
(key == 11'b01100101010) ? 48'b011001010110111010111100000101101111101110101110 :
(key == 11'b01100101011) ? 48'b011001010110011110101001000101101101110000011000 :
(key == 11'b01100101100) ? 48'b011001010110000010011000000101101011110010010000 :
(key == 11'b01100101101) ? 48'b011001010101100110000111100101101001110100010000 :
(key == 11'b01100101110) ? 48'b011001010101001001111000000101100111110110011000 :
(key == 11'b01100101111) ? 48'b011001010100101101101011100101100101111000110010 :
(key == 11'b01100110000) ? 48'b011001010100010001100000000101100011111011010011 :
(key == 11'b01100110001) ? 48'b011001010011110101010101100101100001111110000000 :
(key == 11'b01100110010) ? 48'b011001010011011001001101000101100000000000110111 :
(key == 11'b01100110011) ? 48'b011001010010111101000101100101011110000011111010 :
(key == 11'b01100110100) ? 48'b011001010010100001000000000101011100000111000111 :
(key == 11'b01100110101) ? 48'b011001010010000100111011100101011010001010011111 :
(key == 11'b01100110110) ? 48'b011001010001101000111001000101011000001110000011 :
(key == 11'b01100110111) ? 48'b011001010001001100110111100101010110010001110001 :
(key == 11'b01100111000) ? 48'b011001010000110000110111000101010100010101100111 :
(key == 11'b01100111001) ? 48'b011001010000010100111000000101010010011001101000 :
(key == 11'b01100111010) ? 48'b011001001111111000111011000101010000011101110111 :
(key == 11'b01100111011) ? 48'b011001001111011101000000000101001110100010010010 :
(key == 11'b01100111100) ? 48'b011001001111000001000101100101001100100110110011 :
(key == 11'b01100111101) ? 48'b011001001110100101001101000101001010101011100011 :
(key == 11'b01100111110) ? 48'b011001001110001001010110000101001000110000011011 :
(key == 11'b01100111111) ? 48'b011001001101101101100000000101000110110101011101 :
(key == 11'b01101000000) ? 48'b011001001101010001101100000101000100111010101110 :
(key == 11'b01101000001) ? 48'b011001001100110101111001000101000011000000000110 :
(key == 11'b01101000010) ? 48'b011001001100011010000111100101000001000101101001 :
(key == 11'b01101000011) ? 48'b011001001011111110010111000100111111001011010011 :
(key == 11'b01101000100) ? 48'b011001001011100010101000000100111101010001001100 :
(key == 11'b01101000101) ? 48'b011001001011000110111011000100111011010111001111 :
(key == 11'b01101000110) ? 48'b011001001010101011001111000100111001011101011010 :
(key == 11'b01101000111) ? 48'b011001001010001111100101000100110111100011110011 :
(key == 11'b01101001000) ? 48'b011001001001110011111100100100110101101010010110 :
(key == 11'b01101001001) ? 48'b011001001001011000010100000100110011110000111111 :
(key == 11'b01101001010) ? 48'b011001001000111100101110000100110001110111110100 :
(key == 11'b01101001011) ? 48'b011001001000100001001001000100101111111110110101 :
(key == 11'b01101001100) ? 48'b011001001000000101100110100100101110000110000100 :
(key == 11'b01101001101) ? 48'b011001000111101010000101000100101100001101011010 :
(key == 11'b01101001110) ? 48'b011001000111001110100100000100101010010100110111 :
(key == 11'b01101001111) ? 48'b011001000110110011000101000100101000011100100011 :
(key == 11'b01101010000) ? 48'b011001000110010111100111000100100110100100010110 :
(key == 11'b01101010001) ? 48'b011001000101111100001010100100100100101100010011 :
(key == 11'b01101010010) ? 48'b011001000101100000110000000100100010110100011110 :
(key == 11'b01101010011) ? 48'b011001000101000101010111000100100000111100110010 :
(key == 11'b01101010100) ? 48'b011001000100101001111111000100011111000101001111 :
(key == 11'b01101010101) ? 48'b011001000100001110101000000100011101001101110111 :
(key == 11'b01101010110) ? 48'b011001000011110011010010100100011011010110100110 :
(key == 11'b01101010111) ? 48'b011001000011010111111111000100011001011111100100 :
(key == 11'b01101011000) ? 48'b011001000010111100101100000100010111101000101000 :
(key == 11'b01101011001) ? 48'b011001000010100001011100000100010101110001111011 :
(key == 11'b01101011010) ? 48'b011001000010000110001100000100010011111011010101 :
(key == 11'b01101011011) ? 48'b011001000001101010111110000100010010000100111001 :
(key == 11'b01101011100) ? 48'b011001000001001111110001000100010000001110101000 :
(key == 11'b01101011101) ? 48'b011001000000110100100101000100001110011000011110 :
(key == 11'b01101011110) ? 48'b011001000000011001011011000100001100100010100010 :
(key == 11'b01101011111) ? 48'b011000111111111110010010000100001010101100101101 :
(key == 11'b01101100000) ? 48'b011000111111100011001011100100001000110111000110 :
(key == 11'b01101100001) ? 48'b011000111111001000000101100100000111000001100110 :
(key == 11'b01101100010) ? 48'b011000111110101101000001000100000101001100010001 :
(key == 11'b01101100011) ? 48'b011000111110010001111101000100000011010111000011 :
(key == 11'b01101100100) ? 48'b011000111101110110111100000100000001100010000010 :
(key == 11'b01101100101) ? 48'b011000111101011011111011000011111111101101001001 :
(key == 11'b01101100110) ? 48'b011000111101000000111100100011111101111000011110 :
(key == 11'b01101100111) ? 48'b011000111100100101111111000011111100000011111001 :
(key == 11'b01101101000) ? 48'b011000111100001011000010100011111010001111011111 :
(key == 11'b01101101001) ? 48'b011000111011110000001000000011111000011011010000 :
(key == 11'b01101101010) ? 48'b011000111011010101001110000011110110100111001000 :
(key == 11'b01101101011) ? 48'b011000111010111010010100100011110100110011000110 :
(key == 11'b01101101100) ? 48'b011000111010011111011110000011110010111111010110 :
(key == 11'b01101101101) ? 48'b011000111010000100101001000011110001001011101101 :
(key == 11'b01101101110) ? 48'b011000111001101001110101000011101111011000001110 :
(key == 11'b01101101111) ? 48'b011000111001001111000010000011101101100100111001 :
(key == 11'b01101110000) ? 48'b011000111000110100010000000011101011110001101001 :
(key == 11'b01101110001) ? 48'b011000111000011001100000000011101001111110101001 :
(key == 11'b01101110010) ? 48'b011000110111111110110001100011101000001011110000 :
(key == 11'b01101110011) ? 48'b011000110111100100000011100011100110011000111110 :
(key == 11'b01101110100) ? 48'b011000110111001001011000000011100100100110011010 :
(key == 11'b01101110101) ? 48'b011000110110101110101101000011100010110011111101 :
(key == 11'b01101110110) ? 48'b011000110110010100000011000011100001000001101010 :
(key == 11'b01101110111) ? 48'b011000110101111001011011000011011111001111100001 :
(key == 11'b01101111000) ? 48'b011000110101011110110101000011011101011101100011 :
(key == 11'b01101111001) ? 48'b011000110101000100001111000011011011101011101011 :
(key == 11'b01101111010) ? 48'b011000110100101001101011000011011001111001111110 :
(key == 11'b01101111011) ? 48'b011000110100001111001000000011011000001000011011 :
(key == 11'b01101111100) ? 48'b011000110011110100100111000011010110010111000011 :
(key == 11'b01101111101) ? 48'b011000110011011010000111000011010100100101110100 :
(key == 11'b01101111110) ? 48'b011000110010111111101000000011010010110100101101 :
(key == 11'b01101111111) ? 48'b011000110010100101001010100011010001000011101111 :
(key == 11'b01110000000) ? 48'b011000110010001010101110100011001111010010111100 :
(key == 11'b01110000001) ? 48'b011000110001110000010011000011001101100010010000 :
(key == 11'b01110000010) ? 48'b011000110001010101111001100011001011110001101110 :
(key == 11'b01110000011) ? 48'b011000110000111011100001000011001010000001010110 :
(key == 11'b01110000100) ? 48'b011000110000100001001011000011001000010001001011 :
(key == 11'b01110000101) ? 48'b011000110000000110110110000011000110100001000111 :
(key == 11'b01110000110) ? 48'b011000101111101100100001100011000100110001001010 :
(key == 11'b01110000111) ? 48'b011000101111010010001110100011000011000001011000 :
(key == 11'b01110001000) ? 48'b011000101110110111111100000011000001010001101100 :
(key == 11'b01110001001) ? 48'b011000101110011101101011100010111111100010001010 :
(key == 11'b01110001010) ? 48'b011000101110000011011101000010111101110010110110 :
(key == 11'b01110001011) ? 48'b011000101101101001001111000010111100000011101000 :
(key == 11'b01110001100) ? 48'b011000101101001111000011000010111010010100100101 :
(key == 11'b01110001101) ? 48'b011000101100110100111000000010111000100101101011 :
(key == 11'b01110001110) ? 48'b011000101100011010101110000010110110110110111000 :
(key == 11'b01110001111) ? 48'b011000101100000000100110000010110101001000010000 :
(key == 11'b01110010000) ? 48'b011000101011100110011110000010110011011001101110 :
(key == 11'b01110010001) ? 48'b011000101011001100011000100010110001101011011001 :
(key == 11'b01110010010) ? 48'b011000101010110010010100100010101111111101001110 :
(key == 11'b01110010011) ? 48'b011000101010011000010001000010101110001111001010 :
(key == 11'b01110010100) ? 48'b011000101001111110001111000010101100100001001101 :
(key == 11'b01110010101) ? 48'b011000101001100100001110000010101010110011011010 :
(key == 11'b01110010110) ? 48'b011000101001001010001110000010101001000101110001 :
(key == 11'b01110010111) ? 48'b011000101000110000010000000010100111011000010010 :
(key == 11'b01110011000) ? 48'b011000101000010110010011000010100101101010111001 :
(key == 11'b01110011001) ? 48'b011000100111111100010111000010100011111101101011 :
(key == 11'b01110011010) ? 48'b011000100111100010011110000010100010010000101001 :
(key == 11'b01110011011) ? 48'b011000100111001000100100000010100000100011101011 :
(key == 11'b01110011100) ? 48'b011000100110101110101100000010011110110110110111 :
(key == 11'b01110011101) ? 48'b011000100110010100110110100010011101001010010000 :
(key == 11'b01110011110) ? 48'b011000100101111011000001000010011011011101101101 :
(key == 11'b01110011111) ? 48'b011000100101100001001101000010011001110001010110 :
(key == 11'b01110100000) ? 48'b011000100101000111011010100010011000000101000111 :
(key == 11'b01110100001) ? 48'b011000100100101101101000100010010110011000111110 :
(key == 11'b01110100010) ? 48'b011000100100010011111001000010010100101101000010 :
(key == 11'b01110100011) ? 48'b011000100011111010001010000010010011000001001100 :
(key == 11'b01110100100) ? 48'b011000100011100000011100000010010001010101100000 :
(key == 11'b01110100101) ? 48'b011000100011000110101111100010001111101001111100 :
(key == 11'b01110100110) ? 48'b011000100010101101000100000010001101111110100000 :
(key == 11'b01110100111) ? 48'b011000100010010011011010100010001100010011001111 :
(key == 11'b01110101000) ? 48'b011000100001111001110001100010001010101000000100 :
(key == 11'b01110101001) ? 48'b011000100001100000001011000010001000111101000111 :
(key == 11'b01110101010) ? 48'b011000100001000110100101000010000111010010001111 :
(key == 11'b01110101011) ? 48'b011000100000101101000000000010000101100111100010 :
(key == 11'b01110101100) ? 48'b011000100000010011011100100010000011111100111011 :
(key == 11'b01110101101) ? 48'b011000011111111001111010000010000010010010011110 :
(key == 11'b01110101110) ? 48'b011000011111100000011001000010000000101000000111 :
(key == 11'b01110101111) ? 48'b011000011111000110111001000001111110111101111011 :
(key == 11'b01110110000) ? 48'b011000011110101101011010000001111101010011111000 :
(key == 11'b01110110001) ? 48'b011000011110010011111101000001111011101001111110 :
(key == 11'b01110110010) ? 48'b011000011101111010100001000001111010000000001011 :
(key == 11'b01110110011) ? 48'b011000011101100001000110000001111000010110100010 :
(key == 11'b01110110100) ? 48'b011000011101000111101100000001110110101100111111 :
(key == 11'b01110110101) ? 48'b011000011100101110010100100001110101000011101001 :
(key == 11'b01110110110) ? 48'b011000011100010100111101100001110011011010011010 :
(key == 11'b01110110111) ? 48'b011000011011111011100111000001110001110001010001 :
(key == 11'b01110111000) ? 48'b011000011011100010010010100001110000001000010010 :
(key == 11'b01110111001) ? 48'b011000011011001000111111000001101110011111011100 :
(key == 11'b01110111010) ? 48'b011000011010101111101101000001101100110110101101 :
(key == 11'b01110111011) ? 48'b011000011010010110011011000001101011001110000101 :
(key == 11'b01110111100) ? 48'b011000011001111101001011100001101001100101101001 :
(key == 11'b01110111101) ? 48'b011000011001100011111101100001100111111101010110 :
(key == 11'b01110111110) ? 48'b011000011001001010110000000001100110010101001010 :
(key == 11'b01110111111) ? 48'b011000011000110001100100000001100100101101000101 :
(key == 11'b01111000000) ? 48'b011000011000011000011001000001100011000101001001 :
(key == 11'b01111000001) ? 48'b011000010111111111001110100001100001011101010100 :
(key == 11'b01111000010) ? 48'b011000010111100110000110100001011111110101101011 :
(key == 11'b01111000011) ? 48'b011000010111001100111110100001011110001110000110 :
(key == 11'b01111000100) ? 48'b011000010110110011111001000001011100100110101101 :
(key == 11'b01111000101) ? 48'b011000010110011010110100100001011010111111011101 :
(key == 11'b01111000110) ? 48'b011000010110000001110000000001011001011000010001 :
(key == 11'b01111000111) ? 48'b011000010101101000101101100001010111110001001111 :
(key == 11'b01111001000) ? 48'b011000010101001111101101000001010110001010011001 :
(key == 11'b01111001001) ? 48'b011000010100110110101100100001010100100011100110 :
(key == 11'b01111001010) ? 48'b011000010100011101101101100001010010111100111101 :
(key == 11'b01111001011) ? 48'b011000010100000100110000000001010001010110011101 :
(key == 11'b01111001100) ? 48'b011000010011101011110100000001001111110000000111 :
(key == 11'b01111001101) ? 48'b011000010011010010111001000001001110001001110111 :
(key == 11'b01111001110) ? 48'b011000010010111001111111000001001100100011110000 :
(key == 11'b01111001111) ? 48'b011000010010100001000110000001001010111101110000 :
(key == 11'b01111010000) ? 48'b011000010010001000001110100001001001010111111001 :
(key == 11'b01111010001) ? 48'b011000010001101111011000100001000111110010001100 :
(key == 11'b01111010010) ? 48'b011000010001010110100010100001000110001100100010 :
(key == 11'b01111010011) ? 48'b011000010000111101101111000001000100100111000100 :
(key == 11'b01111010100) ? 48'b011000010000100100111100000001000011000001101101 :
(key == 11'b01111010101) ? 48'b011000010000001100001010000001000001011100011111 :
(key == 11'b01111010110) ? 48'b011000001111110011011001100000111111110111010111 :
(key == 11'b01111010111) ? 48'b011000001111011010101001100000111110010010010110 :
(key == 11'b01111011000) ? 48'b011000001111000001111100100000111100101101100100 :
(key == 11'b01111011001) ? 48'b011000001110101001001111100000111011001000110101 :
(key == 11'b01111011010) ? 48'b011000001110010000100100000000111001100100001111 :
(key == 11'b01111011011) ? 48'b011000001101110111111000100000110111111111101101 :
(key == 11'b01111011100) ? 48'b011000001101011111001111000000110110011011010111 :
(key == 11'b01111011101) ? 48'b011000001101000110100111000000110100110111001000 :
(key == 11'b01111011110) ? 48'b011000001100101110000000000000110011010011000001 :
(key == 11'b01111011111) ? 48'b011000001100010101011010000000110001101111000100 :
(key == 11'b01111100000) ? 48'b011000001011111100110110000000110000001011010000 :
(key == 11'b01111100001) ? 48'b011000001011100100010010000000101110100111100000 :
(key == 11'b01111100010) ? 48'b011000001011001011110000000000101101000011111000 :
(key == 11'b01111100011) ? 48'b011000001010110011001111000000101011100000011010 :
(key == 11'b01111100100) ? 48'b011000001010011010101111000000101001111101000101 :
(key == 11'b01111100101) ? 48'b011000001010000010010000000000101000011001110100 :
(key == 11'b01111100110) ? 48'b011000001001101001110010000000100110110110101011 :
(key == 11'b01111100111) ? 48'b011000001001010001010101000000100101010011101100 :
(key == 11'b01111101000) ? 48'b011000001000111000111001100000100011110000110010 :
(key == 11'b01111101001) ? 48'b011000001000100000011111000000100010001110000010 :
(key == 11'b01111101010) ? 48'b011000001000001000000110100000100000101011011100 :
(key == 11'b01111101011) ? 48'b011000000111101111101110100000011111001000111011 :
(key == 11'b01111101100) ? 48'b011000000111010111011000000000011101100110100100 :
(key == 11'b01111101101) ? 48'b011000000110111111000010000000011100000100010010 :
(key == 11'b01111101110) ? 48'b011000000110100110101110000000011010100010001010 :
(key == 11'b01111101111) ? 48'b011000000110001110011010100000011001000000001000 :
(key == 11'b01111110000) ? 48'b011000000101110110001000100000010111011110001111 :
(key == 11'b01111110001) ? 48'b011000000101011101110111000000010101111100011100 :
(key == 11'b01111110010) ? 48'b011000000101000101100111100000010100011010110010 :
(key == 11'b01111110011) ? 48'b011000000100101101011000100000010010111001001111 :
(key == 11'b01111110100) ? 48'b011000000100010101001011000000010001010111110100 :
(key == 11'b01111110101) ? 48'b011000000011111100111110000000001111110110100000 :
(key == 11'b01111110110) ? 48'b011000000011100100110011000000001110010101010100 :
(key == 11'b01111110111) ? 48'b011000000011001100101001000000001100110100010010 :
(key == 11'b01111111000) ? 48'b011000000010110100100000000000001011010011010110 :
(key == 11'b01111111001) ? 48'b011000000010011100011000000000001001110010100000 :
(key == 11'b01111111010) ? 48'b011000000010000100010001000000001000010001110011 :
(key == 11'b01111111011) ? 48'b011000000001101100001011000000000110110001001011 :
(key == 11'b01111111100) ? 48'b011000000001010100000111100000000101010000110000 :
(key == 11'b01111111101) ? 48'b011000000000111100000100000000000011110000011000 :
(key == 11'b01111111110) ? 48'b011000000000100100000001100000000010010000001001 :
(key == 11'b01111111111) ? 48'b011000000000001100000001000000000000110000000011 :
(key == 11'b10000000000) ? 48'b101111111111010000000010011111111101000000001100 :
(key == 11'b10000000001) ? 48'b101111111101110000001011011111110111000001001000 :
(key == 11'b10000000010) ? 48'b101111111100010000011101011111110001000011000000 :
(key == 11'b10000000011) ? 48'b101111111010110000111000011111101011000101110011 :
(key == 11'b10000000100) ? 48'b101111111001010001011100011111100101001001100010 :
(key == 11'b10000000101) ? 48'b101111110111110010001000011111011111001110001010 :
(key == 11'b10000000110) ? 48'b101111110110010010111110011111011001010011110000 :
(key == 11'b10000000111) ? 48'b101111110100110011111110011111010011011010010001 :
(key == 11'b10000001000) ? 48'b101111110011010101000100011111001101100001100111 :
(key == 11'b10000001001) ? 48'b101111110001110110010101011111000111101001111110 :
(key == 11'b10000001010) ? 48'b101111110000010111101110011111000001110011001011 :
(key == 11'b10000001011) ? 48'b101111101110111001001110011110111011111101001111 :
(key == 11'b10000001100) ? 48'b101111101101011010111010011110110110001000010011 :
(key == 11'b10000001101) ? 48'b101111101011111100101101011110110000010100010000 :
(key == 11'b10000001110) ? 48'b101111101010011110101000011110101010100001000000 :
(key == 11'b10000001111) ? 48'b101111101001000000101100011110100100101110101100 :
(key == 11'b10000010000) ? 48'b101111100111100010111010011110011110111101010111 :
(key == 11'b10000010001) ? 48'b101111100110000101010000011110011001001100110111 :
(key == 11'b10000010010) ? 48'b101111100100100111101111011110010011011101001101 :
(key == 11'b10000010011) ? 48'b101111100011001010010110011110001101101110011110 :
(key == 11'b10000010100) ? 48'b101111100001101101000110011110001000000000100101 :
(key == 11'b10000010101) ? 48'b101111100000001111111110011110000010010011100110 :
(key == 11'b10000010110) ? 48'b101111011110110010111110011101111100100111011011 :
(key == 11'b10000010111) ? 48'b101111011101010110000111011101110110111100001001 :
(key == 11'b10000011000) ? 48'b101111011011111001011001011101110001010001110000 :
(key == 11'b10000011001) ? 48'b101111011010011100110100011101101011101000010001 :
(key == 11'b10000011010) ? 48'b101111011001000000010111011101100101111111101000 :
(key == 11'b10000011011) ? 48'b101111010111100100000010011101100000010111110010 :
(key == 11'b10000011100) ? 48'b101111010110000111110101011101011010110000110011 :
(key == 11'b10000011101) ? 48'b101111010100101011110001011101010101001010101100 :
(key == 11'b10000011110) ? 48'b101111010011001111110110011101001111100101011110 :
(key == 11'b10000011111) ? 48'b101111010001110100000010011101001010000001000010 :
(key == 11'b10000100000) ? 48'b101111010000011000011000011101000100011101011111 :
(key == 11'b10000100001) ? 48'b101111001110111100110101011100111110111010101111 :
(key == 11'b10000100010) ? 48'b101111001101100001011011011100111001011000110111 :
(key == 11'b10000100011) ? 48'b101111001100000110001010011100110011110111110111 :
(key == 11'b10000100100) ? 48'b101111001010101011000000011100101110010111101010 :
(key == 11'b10000100101) ? 48'b101111001001001111111110011100101000111000001110 :
(key == 11'b10000100110) ? 48'b101111000111110101000110011100100011011001101011 :
(key == 11'b10000100111) ? 48'b101111000110011010010100011100011101111011111001 :
(key == 11'b10000101000) ? 48'b101111000100111111101011011100011000011110111101 :
(key == 11'b10000101001) ? 48'b101111000011100101001010011100010011000010111000 :
(key == 11'b10000101010) ? 48'b101111000010001010110010011100001101100111100100 :
(key == 11'b10000101011) ? 48'b101111000000110000100000011100001000001101000011 :
(key == 11'b10000101100) ? 48'b101110111111010110011001011100000010110011011011 :
(key == 11'b10000101101) ? 48'b101110111101111100011001011011111101011010100101 :
(key == 11'b10000101110) ? 48'b101110111100100010100001011011111000000010100011 :
(key == 11'b10000101111) ? 48'b101110111011001000110001011011110010101011010010 :
(key == 11'b10000110000) ? 48'b101110111001101111001001011011101101010100110110 :
(key == 11'b10000110001) ? 48'b101110111000010101101000011011100111111111001010 :
(key == 11'b10000110010) ? 48'b101110110110111100010001011011100010101010010101 :
(key == 11'b10000110011) ? 48'b101110110101100011000001011011011101010110010001 :
(key == 11'b10000110100) ? 48'b101110110100001001111000011011011000000010111110 :
(key == 11'b10000110101) ? 48'b101110110010110000111001011011010010110000100001 :
(key == 11'b10000110110) ? 48'b101110110001011000000001011011001101011110110100 :
(key == 11'b10000110111) ? 48'b101110101111111111010000011011001000001101110110 :
(key == 11'b10000111000) ? 48'b101110101110100110101000011011000010111101101110 :
(key == 11'b10000111001) ? 48'b101110101101001110001000011010111101101110011000 :
(key == 11'b10000111010) ? 48'b101110101011110101101111011010111000011111110011 :
(key == 11'b10000111011) ? 48'b101110101010011101011110011010110011010001111110 :
(key == 11'b10000111100) ? 48'b101110101001000101010100011010101110000100111001 :
(key == 11'b10000111101) ? 48'b101110100111101101010100011010101000111000101010 :
(key == 11'b10000111110) ? 48'b101110100110010101011010011010100011101101000111 :
(key == 11'b10000111111) ? 48'b101110100100111101101001011010011110100010011000 :
(key == 11'b10001000000) ? 48'b101110100011100110000000011010011001011000011010 :
(key == 11'b10001000001) ? 48'b101110100010001110011101011010010100001111001010 :
(key == 11'b10001000010) ? 48'b101110100000110111000010011010001111000110101001 :
(key == 11'b10001000011) ? 48'b101110011111011111110000011010001001111110111101 :
(key == 11'b10001000100) ? 48'b101110011110001000100100011010000100110111111011 :
(key == 11'b10001000101) ? 48'b101110011100110001100000011001111111110001101011 :
(key == 11'b10001000110) ? 48'b101110011011011010100100011001111010101100001010 :
(key == 11'b10001000111) ? 48'b101110011010000011110000011001110101100111011011 :
(key == 11'b10001001000) ? 48'b101110011000101101000100011001110000100011011011 :
(key == 11'b10001001001) ? 48'b101110010111010110011111011001101011100000001101 :
(key == 11'b10001001010) ? 48'b101110010110000000000010011001100110011101101011 :
(key == 11'b10001001011) ? 48'b101110010100101001101011011001100001011011110100 :
(key == 11'b10001001100) ? 48'b101110010011010011011100011001011100011010101111 :
(key == 11'b10001001101) ? 48'b101110010001111101010110011001010111011010011100 :
(key == 11'b10001001110) ? 48'b101110010000100111010111011001010010011010110100 :
(key == 11'b10001001111) ? 48'b101110001111010001011111011001001101011011111011 :
(key == 11'b10001010000) ? 48'b101110001101111011101111011001001000011101110010 :
(key == 11'b10001010001) ? 48'b101110001100100110000110011001000011100000010101 :
(key == 11'b10001010010) ? 48'b101110001011010000100100011000111110100011100110 :
(key == 11'b10001010011) ? 48'b101110001001111011001010011000111001100111100011 :
(key == 11'b10001010100) ? 48'b101110001000100101110111011000110100101100010000 :
(key == 11'b10001010101) ? 48'b101110000111010000101100011000101111110001101001 :
(key == 11'b10001010110) ? 48'b101110000101111011101000011000101010110111110010 :
(key == 11'b10001010111) ? 48'b101110000100100110101011011000100101111110100110 :
(key == 11'b10001011000) ? 48'b101110000011010001110110011000100001000110000111 :
(key == 11'b10001011001) ? 48'b101110000001111101001000011000011100001110010100 :
(key == 11'b10001011010) ? 48'b101110000000101000100000011000010111010111001110 :
(key == 11'b10001011011) ? 48'b101101111111010100000010011000010010100000111000 :
(key == 11'b10001011100) ? 48'b101101111101111111101010011000001101101011001100 :
(key == 11'b10001011101) ? 48'b101101111100101011011000011000001000110110001100 :
(key == 11'b10001011110) ? 48'b101101111011010111001111011000000100000001111000 :
(key == 11'b10001011111) ? 48'b101101111010000011001100010111111111001110010001 :
(key == 11'b10001100000) ? 48'b101101111000101111010001010111111010011011010101 :
(key == 11'b10001100001) ? 48'b101101110111011011011101010111110101101001000110 :
(key == 11'b10001100010) ? 48'b101101110110000111110000010111110000110111100011 :
(key == 11'b10001100011) ? 48'b101101110100110100001011010111101100000110101010 :
(key == 11'b10001100100) ? 48'b101101110011100000101100010111100111010110011110 :
(key == 11'b10001100101) ? 48'b101101110010001101010101010111100010100110111100 :
(key == 11'b10001100110) ? 48'b101101110000111010000100010111011101111000000100 :
(key == 11'b10001100111) ? 48'b101101101111100110111011010111011001001001111000 :
(key == 11'b10001101000) ? 48'b101101101110010011111000010111010100011100010110 :
(key == 11'b10001101001) ? 48'b101101101101000000111110010111001111101111100100 :
(key == 11'b10001101010) ? 48'b101101101011101110001010010111001011000011011000 :
(key == 11'b10001101011) ? 48'b101101101010011011011100010111000110010111110100 :
(key == 11'b10001101100) ? 48'b101101101001001000110110010111000001101100111110 :
(key == 11'b10001101101) ? 48'b101101100111110110011000010110111101000010110011 :
(key == 11'b10001101110) ? 48'b101101100110100100000000010110111000011001001111 :
(key == 11'b10001101111) ? 48'b101101100101010001101110010110110011110000010110 :
(key == 11'b10001110000) ? 48'b101101100011111111100101010110101111001000001010 :
(key == 11'b10001110001) ? 48'b101101100010101101100001010110101010100000100001 :
(key == 11'b10001110010) ? 48'b101101100001011011100100010110100101111001100011 :
(key == 11'b10001110011) ? 48'b101101100000001001110000010110100001010011010100 :
(key == 11'b10001110100) ? 48'b101101011110111000000001010110011100101101101011 :
(key == 11'b10001110101) ? 48'b101101011101100110011000010110011000001000101000 :
(key == 11'b10001110110) ? 48'b101101011100010100111000010110010011100100010000 :
(key == 11'b10001110111) ? 48'b101101011011000011011110010110001111000000100100 :
(key == 11'b10001111000) ? 48'b101101011001110010001010010110001010011101011101 :
(key == 11'b10001111001) ? 48'b101101011000100000111110010110000101111011000001 :
(key == 11'b10001111010) ? 48'b101101010111001111111000010110000001011001001011 :
(key == 11'b10001111011) ? 48'b101101010101111110111010010101111100111000000000 :
(key == 11'b10001111100) ? 48'b101101010100101110000011010101111000010111100000 :
(key == 11'b10001111101) ? 48'b101101010011011101010001010101110011110111100011 :
(key == 11'b10001111110) ? 48'b101101010010001100100111010101101111011000010000 :
(key == 11'b10001111111) ? 48'b101101010000111100000100010101101010111001100110 :
(key == 11'b10010000000) ? 48'b101101001111101011101000010101100110011011100110 :
(key == 11'b10010000001) ? 48'b101101001110011011010000010101100001111110000110 :
(key == 11'b10010000010) ? 48'b101101001101001011000000010101011101100001010000 :
(key == 11'b10010000011) ? 48'b101101001011111010111000010101011001000101000100 :
(key == 11'b10010000100) ? 48'b101101001010101010110101010101010100101001011110 :
(key == 11'b10010000101) ? 48'b101101001001011010111010010101010000001110100010 :
(key == 11'b10010000110) ? 48'b101101001000001011000100010101001011110100001000 :
(key == 11'b10010000111) ? 48'b101101000110111011010110010101000111011010011000 :
(key == 11'b10010001000) ? 48'b101101000101101011101110010101000011000001010000 :
(key == 11'b10010001001) ? 48'b101101000100011100001110010100111110101000101111 :
(key == 11'b10010001010) ? 48'b101101000011001100110010010100111010010000110000 :
(key == 11'b10010001011) ? 48'b101101000001111101011110010100110101111001011010 :
(key == 11'b10010001100) ? 48'b101101000000101110010001010100110001100010101100 :
(key == 11'b10010001101) ? 48'b101100111111011111001001010100101101001100100000 :
(key == 11'b10010001110) ? 48'b101100111110010000001000010100101000110110111101 :
(key == 11'b10010001111) ? 48'b101100111101000001010000010100100100100010000100 :
(key == 11'b10010010000) ? 48'b101100111011110010011011010100100000001101101010 :
(key == 11'b10010010001) ? 48'b101100111010100011101110010100011011111001111000 :
(key == 11'b10010010010) ? 48'b101100111001010101001000010100010111100110101111 :
(key == 11'b10010010011) ? 48'b101100111000000110101000010100010011010100001000 :
(key == 11'b10010010100) ? 48'b101100110110111000001110010100001111000010001001 :
(key == 11'b10010010101) ? 48'b101100110101101001111010010100001010110000101101 :
(key == 11'b10010010110) ? 48'b101100110100011011101101010100000110011111110101 :
(key == 11'b10010010111) ? 48'b101100110011001101100111010100000010001111100110 :
(key == 11'b10010011000) ? 48'b101100110001111111100110010011111101111111111001 :
(key == 11'b10010011001) ? 48'b101100110000110001101100010011111001110000110001 :
(key == 11'b10010011010) ? 48'b101100101111100011111001010011110101100010010000 :
(key == 11'b10010011011) ? 48'b101100101110010110001100010011110001010100010101 :
(key == 11'b10010011100) ? 48'b101100101101001000100110010011101101000110111110 :
(key == 11'b10010011101) ? 48'b101100101011111011000110010011101000111010001001 :
(key == 11'b10010011110) ? 48'b101100101010101101101011010011100100101101111000 :
(key == 11'b10010011111) ? 48'b101100101001100000010110010011100000100010001010 :
(key == 11'b10010100000) ? 48'b101100101000010011001010010011011100010111000110 :
(key == 11'b10010100001) ? 48'b101100100111000110000010010011011000001100100100 :
(key == 11'b10010100010) ? 48'b101100100101111001000001010011010100000010100010 :
(key == 11'b10010100011) ? 48'b101100100100101100000110010011001111111001000110 :
(key == 11'b10010100100) ? 48'b101100100011011111010001010011001011110000001101 :
(key == 11'b10010100101) ? 48'b101100100010010010100010010011000111100111111010 :
(key == 11'b10010100110) ? 48'b101100100001000101111010010011000011100000000110 :
(key == 11'b10010100111) ? 48'b101100011111111001011000010010111111011000111100 :
(key == 11'b10010101000) ? 48'b101100011110101100111100010010111011010010010000 :
(key == 11'b10010101001) ? 48'b101100011101100000100110010010110111001100001000 :
(key == 11'b10010101010) ? 48'b101100011100010100010110010010110011000110100101 :
(key == 11'b10010101011) ? 48'b101100011011001000001100010010101111000001100100 :
(key == 11'b10010101100) ? 48'b101100011001111100001001010010101010111101000110 :
(key == 11'b10010101101) ? 48'b101100011000110000001100010010100110111001001011 :
(key == 11'b10010101110) ? 48'b101100010111100100010100010010100010110101110010 :
(key == 11'b10010101111) ? 48'b101100010110011000100010010010011110110010111100 :
(key == 11'b10010110000) ? 48'b101100010101001100111000010010011010110000101100 :
(key == 11'b10010110001) ? 48'b101100010100000001010011010010010110101110111010 :
(key == 11'b10010110010) ? 48'b101100010010110101110100010010010010101101101010 :
(key == 11'b10010110011) ? 48'b101100010001101010011010010010001110101100111100 :
(key == 11'b10010110100) ? 48'b101100010000011111001000010010001010101100110100 :
(key == 11'b10010110101) ? 48'b101100001111010011111010010010000110101101001011 :
(key == 11'b10010110110) ? 48'b101100001110001000110011010010000010101110000011 :
(key == 11'b10010110111) ? 48'b101100001100111101110011010001111110101111100010 :
(key == 11'b10010111000) ? 48'b101100001011110010111000010001111010110001011110 :
(key == 11'b10010111001) ? 48'b101100001010101000000011010001110110110011111110 :
(key == 11'b10010111010) ? 48'b101100001001011101010010010001110010110110111010 :
(key == 11'b10010111011) ? 48'b101100001000010010101001010001101110111010011100 :
(key == 11'b10010111100) ? 48'b101100000111001000000111010001101010111110100011 :
(key == 11'b10010111101) ? 48'b101100000101111101101010010001100111000011000111 :
(key == 11'b10010111110) ? 48'b101100000100110011010001010001100011001000001010 :
(key == 11'b10010111111) ? 48'b101100000011101000111111010001011111001101101110 :
(key == 11'b10011000000) ? 48'b101100000010011110110100010001011011010011110111 :
(key == 11'b10011000001) ? 48'b101100000001010100101101010001010111011010011110 :
(key == 11'b10011000010) ? 48'b101100000000001010101101010001010011100001100111 :
(key == 11'b10011000011) ? 48'b101011111111000000110100010001001111101001010011 :
(key == 11'b10011000100) ? 48'b101011111101110110111110010001001011110001011011 :
(key == 11'b10011000101) ? 48'b101011111100101101010000010001000111111010000101 :
(key == 11'b10011000110) ? 48'b101011111011100011100110010001000100000011001111 :
(key == 11'b10011000111) ? 48'b101011111010011010000100010001000000001100111100 :
(key == 11'b10011001000) ? 48'b101011111001010000100110010000111100010111001000 :
(key == 11'b10011001001) ? 48'b101011111000000111001110010000111000100001110000 :
(key == 11'b10011001010) ? 48'b101011110110111101111100010000110100101100111100 :
(key == 11'b10011001011) ? 48'b101011110101110100110000010000110000111000100110 :
(key == 11'b10011001100) ? 48'b101011110100101011101010010000101101000100110011 :
(key == 11'b10011001101) ? 48'b101011110011100010101001010000101001010001011100 :
(key == 11'b10011001110) ? 48'b101011110010011001101110010000100101011110100110 :
(key == 11'b10011001111) ? 48'b101011110001010000111001010000100001101100010011 :
(key == 11'b10011010000) ? 48'b101011110000001000001001010000011101111010011011 :
(key == 11'b10011010001) ? 48'b101011101110111111011110010000011010001001000010 :
(key == 11'b10011010010) ? 48'b101011101101110110111010010000010110011000001010 :
(key == 11'b10011010011) ? 48'b101011101100101110011100010000010010100111110010 :
(key == 11'b10011010100) ? 48'b101011101011100110000100010000001110110111111100 :
(key == 11'b10011010101) ? 48'b101011101010011101110000010000001011001000100001 :
(key == 11'b10011010110) ? 48'b101011101001010101100001010000000111011001100010 :
(key == 11'b10011010111) ? 48'b101011101000001101011000010000000011101011000010 :
(key == 11'b10011011000) ? 48'b101011100111000101010110001111111111111101001000 :
(key == 11'b10011011001) ? 48'b101011100101111101011010001111111100001111101000 :
(key == 11'b10011011010) ? 48'b101011100100110101100001001111111000100010100101 :
(key == 11'b10011011011) ? 48'b101011100011101101101110001111110100110110000001 :
(key == 11'b10011011100) ? 48'b101011100010100110000011001111110001001001111111 :
(key == 11'b10011011101) ? 48'b101011100001011110011100001111101101011110011000 :
(key == 11'b10011011110) ? 48'b101011100000010110111011001111101001110011010100 :
(key == 11'b10011011111) ? 48'b101011011111001111011111001111100110001000101010 :
(key == 11'b10011100000) ? 48'b101011011110001000001000001111100010011110011110 :
(key == 11'b10011100001) ? 48'b101011011101000000111000001111011110110100110001 :
(key == 11'b10011100010) ? 48'b101011011011111001101011001111011011001011100000 :
(key == 11'b10011100011) ? 48'b101011011010110010100101001111010111100010101101 :
(key == 11'b10011100100) ? 48'b101011011001101011100101001111010011111010011010 :
(key == 11'b10011100101) ? 48'b101011011000100100101010001111010000010010100111 :
(key == 11'b10011100110) ? 48'b101011010111011101110100001111001100101011001100 :
(key == 11'b10011100111) ? 48'b101011010110010111000100001111001001000100010000 :
(key == 11'b10011101000) ? 48'b101011010101010000011001001111000101011101110100 :
(key == 11'b10011101001) ? 48'b101011010100001001110011001111000001110111110001 :
(key == 11'b10011101010) ? 48'b101011010011000011010011001110111110010010001110 :
(key == 11'b10011101011) ? 48'b101011010001111100111000001110111010101101000110 :
(key == 11'b10011101100) ? 48'b101011010000110110100011001110110111001000011110 :
(key == 11'b10011101101) ? 48'b101011001111110000010010001110110011100100010010 :
(key == 11'b10011101110) ? 48'b101011001110101010001000001110110000000000100100 :
(key == 11'b10011101111) ? 48'b101011001101100100000011001110101100011101010011 :
(key == 11'b10011110000) ? 48'b101011001100011110000100001110101000111010011110 :
(key == 11'b10011110001) ? 48'b101011001011011000001000001110100101011000000100 :
(key == 11'b10011110010) ? 48'b101011001010010010010011001110100001110110001000 :
(key == 11'b10011110011) ? 48'b101011001001001100100011001110011110010100101000 :
(key == 11'b10011110100) ? 48'b101011001000000110111000001110011010110011100100 :
(key == 11'b10011110101) ? 48'b101011000111000001010010001110010111010010111100 :
(key == 11'b10011110110) ? 48'b101011000101111011110010001110010011110010110100 :
(key == 11'b10011110111) ? 48'b101011000100110110010111001110010000010011000100 :
(key == 11'b10011111000) ? 48'b101011000011110001000001001110001100110011110010 :
(key == 11'b10011111001) ? 48'b101011000010101011110000001110001001010100111100 :
(key == 11'b10011111010) ? 48'b101011000001100110100100001110000101110110011111 :
(key == 11'b10011111011) ? 48'b101011000000100001011110001110000010011000100001 :
(key == 11'b10011111100) ? 48'b101010111111011100011110001101111110111011000000 :
(key == 11'b10011111101) ? 48'b101010111110010111100010001101111011011101110111 :
(key == 11'b10011111110) ? 48'b101010111101010010101011001101111000000001001101 :
(key == 11'b10011111111) ? 48'b101010111100001101111010001101110100100100111100 :
(key == 11'b10100000000) ? 48'b101010111011001001001101001101110001001001001000 :
(key == 11'b10100000001) ? 48'b101010111010000100100110001101101101101101110001 :
(key == 11'b10100000010) ? 48'b101010111001000000000100001101101010010010110011 :
(key == 11'b10100000011) ? 48'b101010110111111011101000001101100110111000010010 :
(key == 11'b10100000100) ? 48'b101010110110110111010000001101100011011110001010 :
(key == 11'b10100000101) ? 48'b101010110101110010111100001101100000000100011100 :
(key == 11'b10100000110) ? 48'b101010110100101110110000001101011100101011001110 :
(key == 11'b10100000111) ? 48'b101010110011101010100111001101011001010010011000 :
(key == 11'b10100001000) ? 48'b101010110010100110100100001101010101111010000000 :
(key == 11'b10100001001) ? 48'b101010110001100010100110001101010010100010000010 :
(key == 11'b10100001010) ? 48'b101010110000011110101101001101001111001010011100 :
(key == 11'b10100001011) ? 48'b101010101111011010111000001101001011110011001111 :
(key == 11'b10100001100) ? 48'b101010101110010111001001001101001000011100100000 :
(key == 11'b10100001101) ? 48'b101010101101010011011110001101000101000110001010 :
(key == 11'b10100001110) ? 48'b101010101100001111111010001101000001110000010000 :
(key == 11'b10100001111) ? 48'b101010101011001100011010001100111110011010110001 :
(key == 11'b10100010000) ? 48'b101010101010001000111110001100111011000101101010 :
(key == 11'b10100010001) ? 48'b101010101001000101101000001100110111110000111110 :
(key == 11'b10100010010) ? 48'b101010101000000010010111001100110100011100101101 :
(key == 11'b10100010011) ? 48'b101010100110111111001100001100110001001000110111 :
(key == 11'b10100010100) ? 48'b101010100101111100000100001100101101110101010111 :
(key == 11'b10100010101) ? 48'b101010100100111001000010001100101010100010010100 :
(key == 11'b10100010110) ? 48'b101010100011110110000100001100100111001111101011 :
(key == 11'b10100010111) ? 48'b101010100010110011001100001100100011111101011100 :
(key == 11'b10100011000) ? 48'b101010100001110000011000001100100000101011100110 :
(key == 11'b10100011001) ? 48'b101010100000101101101010001100011101011010001010 :
(key == 11'b10100011010) ? 48'b101010011111101011000000001100011010001001001000 :
(key == 11'b10100011011) ? 48'b101010011110101000011100001100010110111000100000 :
(key == 11'b10100011100) ? 48'b101010011101100101111100001100010011101000010010 :
(key == 11'b10100011101) ? 48'b101010011100100011100000001100010000011000011001 :
(key == 11'b10100011110) ? 48'b101010011011100001001010001100001101001000111110 :
(key == 11'b10100011111) ? 48'b101010011010011110111000001100001001111001111001 :
(key == 11'b10100100000) ? 48'b101010011001011100101100001100000110101011010000 :
(key == 11'b10100100001) ? 48'b101010011000011010100101001100000011011101000000 :
(key == 11'b10100100010) ? 48'b101010010111011000100010001100000000001111000111 :
(key == 11'b10100100011) ? 48'b101010010110010110100100001011111101000001101001 :
(key == 11'b10100100100) ? 48'b101010010101010100101011001011111001110100100011 :
(key == 11'b10100100101) ? 48'b101010010100010010110111001011110110100111111000 :
(key == 11'b10100100110) ? 48'b101010010011010001001000001011110011011011100100 :
(key == 11'b10100100111) ? 48'b101010010010001111011100001011110000001111101000 :
(key == 11'b10100101000) ? 48'b101010010001001101110111001011101101000100000110 :
(key == 11'b10100101001) ? 48'b101010010000001100010110001011101001111000111100 :
(key == 11'b10100101010) ? 48'b101010001111001010111010001011100110101110001100 :
(key == 11'b10100101011) ? 48'b101010001110001001100001001011100011100011110010 :
(key == 11'b10100101100) ? 48'b101010001101001000001110001011100000011001101111 :
(key == 11'b10100101101) ? 48'b101010001100000110111111001011011101010000000110 :
(key == 11'b10100101110) ? 48'b101010001011000101110110001011011010000110110111 :
(key == 11'b10100101111) ? 48'b101010001010000100110001001011010110111110000000 :
(key == 11'b10100110000) ? 48'b101010001001000011110010001011010011110101100011 :
(key == 11'b10100110001) ? 48'b101010001000000010110110001011010000101101011011 :
(key == 11'b10100110010) ? 48'b101010000111000001111111001011001101100101101100 :
(key == 11'b10100110011) ? 48'b101010000110000001001110001011001010011110011000 :
(key == 11'b10100110100) ? 48'b101010000101000000100000001011000111010111010110 :
(key == 11'b10100110101) ? 48'b101010000011111111110111001011000100010000101110 :
(key == 11'b10100110110) ? 48'b101010000010111111010011001011000001001010100000 :
(key == 11'b10100110111) ? 48'b101010000001111110110011001010111110000100100110 :
(key == 11'b10100111000) ? 48'b101010000000111110011001001010111010111111001001 :
(key == 11'b10100111001) ? 48'b101001111111111110000011001010110111111010000000 :
(key == 11'b10100111010) ? 48'b101001111110111101110001001010110100110101001111 :
(key == 11'b10100111011) ? 48'b101001111101111101100100001010110001110000110111 :
(key == 11'b10100111100) ? 48'b101001111100111101011100001010101110101100110100 :
(key == 11'b10100111101) ? 48'b101001111011111101011000001010101011101001001000 :
(key == 11'b10100111110) ? 48'b101001111010111101011000001010101000100101110110 :
(key == 11'b10100111111) ? 48'b101001111001111101011110001010100101100010111010 :
(key == 11'b10101000000) ? 48'b101001111000111101101000001010100010100000010101 :
(key == 11'b10101000001) ? 48'b101001110111111101110110001010011111011110001000 :
(key == 11'b10101000010) ? 48'b101001110110111110001010001010011100011100010001 :
(key == 11'b10101000011) ? 48'b101001110101111110100001001010011001011010110001 :
(key == 11'b10101000100) ? 48'b101001110100111110111101001010010110011001101000 :
(key == 11'b10101000101) ? 48'b101001110011111111011110001010010011011000110110 :
(key == 11'b10101000110) ? 48'b101001110011000000000011001010010000011000011110 :
(key == 11'b10101000111) ? 48'b101001110010000000101101001010001101011000011000 :
(key == 11'b10101001000) ? 48'b101001110001000001011011001010001010011000101011 :
(key == 11'b10101001001) ? 48'b101001110000000010001110001010000111011001010110 :
(key == 11'b10101001010) ? 48'b101001101111000011000101001010000100011010010101 :
(key == 11'b10101001011) ? 48'b101001101110000100000000001010000001011011101100 :
(key == 11'b10101001100) ? 48'b101001101101000101000000001001111110011101011001 :
(key == 11'b10101001101) ? 48'b101001101100000110000101001001111011011111011100 :
(key == 11'b10101001110) ? 48'b101001101011000111001110001001111000100001110110 :
(key == 11'b10101001111) ? 48'b101001101010001000011100001001110101100100100110 :
(key == 11'b10101010000) ? 48'b101001101001001001101110001001110010100111101101 :
(key == 11'b10101010001) ? 48'b101001101000001011000100001001101111101011001010 :
(key == 11'b10101010010) ? 48'b101001100111001100011110001001101100101110111011 :
(key == 11'b10101010011) ? 48'b101001100110001101111101001001101001110011000011 :
(key == 11'b10101010100) ? 48'b101001100101001111100001001001100110110111100100 :
(key == 11'b10101010101) ? 48'b101001100100010001001001001001100011111100011000 :
(key == 11'b10101010110) ? 48'b101001100011010010110101001001100001000001100010 :
(key == 11'b10101010111) ? 48'b101001100010010100100110001001011110000111000101 :
(key == 11'b10101011000) ? 48'b101001100001010110011011001001011011001100111010 :
(key == 11'b10101011001) ? 48'b101001100000011000010100001001011000010011000101 :
(key == 11'b10101011010) ? 48'b101001011111011010010010001001010101011001101000 :
(key == 11'b10101011011) ? 48'b101001011110011100010100001001010010100000011111 :
(key == 11'b10101011100) ? 48'b101001011101011110011010001001001111100111101010 :
(key == 11'b10101011101) ? 48'b101001011100100000100101001001001100101111001110 :
(key == 11'b10101011110) ? 48'b101001011011100010110100001001001001110111000111 :
(key == 11'b10101011111) ? 48'b101001011010100101000111001001000110111111010010 :
(key == 11'b10101100000) ? 48'b101001011001100111100000001001000100000111110111 :
(key == 11'b10101100001) ? 48'b101001011000101001111011001001000001010000101110 :
(key == 11'b10101100010) ? 48'b101001010111101100011100001000111110011001111100 :
(key == 11'b10101100011) ? 48'b101001010110101111000001001000111011100011100001 :
(key == 11'b10101100100) ? 48'b101001010101110001101001001000111000101101010111 :
(key == 11'b10101100101) ? 48'b101001010100110100010110001000110101110111100011 :
(key == 11'b10101100110) ? 48'b101001010011110111000110001000110011000010000010 :
(key == 11'b10101100111) ? 48'b101001010010111001111100001000110000001100111001 :
(key == 11'b10101101000) ? 48'b101001010001111100110110001000101101011000000110 :
(key == 11'b10101101001) ? 48'b101001010000111111110100001000101010100011100110 :
(key == 11'b10101101010) ? 48'b101001010000000010110111001000100111101111011101 :
(key == 11'b10101101011) ? 48'b101001001111000101111101001000100100111011100110 :
(key == 11'b10101101100) ? 48'b101001001110001001001000001000100010001000000101 :
(key == 11'b10101101101) ? 48'b101001001101001100010111001000011111010100111010 :
(key == 11'b10101101110) ? 48'b101001001100001111101010001000011100100010000001 :
(key == 11'b10101101111) ? 48'b101001001011010011000001001000011001101111011101 :
(key == 11'b10101110000) ? 48'b101001001010010110011101001000010110111101001111 :
(key == 11'b10101110001) ? 48'b101001001001011001111101001000010100001011010101 :
(key == 11'b10101110010) ? 48'b101001001000011101100001001000010001011001110000 :
(key == 11'b10101110011) ? 48'b101001000111100001001001001000001110101000011111 :
(key == 11'b10101110100) ? 48'b101001000110100100110100001000001011110111011111 :
(key == 11'b10101110101) ? 48'b101001000101101000100100001000001001000110110110 :
(key == 11'b10101110110) ? 48'b101001000100101100011001001000000110010110100010 :
(key == 11'b10101110111) ? 48'b101001000011110000010010001000000011100110100001 :
(key == 11'b10101111000) ? 48'b101001000010110100001110001000000000110110110110 :
(key == 11'b10101111001) ? 48'b101001000001111000001111000111111110000111011101 :
(key == 11'b10101111010) ? 48'b101001000000111100010100000111111011011000011010 :
(key == 11'b10101111011) ? 48'b101001000000000000011101000111111000101001100111 :
(key == 11'b10101111100) ? 48'b101000111111000100101010000111110101111011001001 :
(key == 11'b10101111101) ? 48'b101000111110001000111100000111110011001101000011 :
(key == 11'b10101111110) ? 48'b101000111101001101010000000111110000011111001101 :
(key == 11'b10101111111) ? 48'b101000111100010001101010000111101101110001101101 :
(key == 11'b10110000000) ? 48'b101000111011010110000111000111101011000100011111 :
(key == 11'b10110000001) ? 48'b101000111010011010101001000111101000010111100110 :
(key == 11'b10110000010) ? 48'b101000111001011111001110000111100101101011000000 :
(key == 11'b10110000011) ? 48'b101000111000100011111000000111100010111110101101 :
(key == 11'b10110000100) ? 48'b101000110111101000100110000111100000010010101110 :
(key == 11'b10110000101) ? 48'b101000110110101101010111000111011101100111000010 :
(key == 11'b10110000110) ? 48'b101000110101110010001100000111011010111011101001 :
(key == 11'b10110000111) ? 48'b101000110100110111000110000111011000010000100100 :
(key == 11'b10110001000) ? 48'b101000110011111100000100000111010101100101110010 :
(key == 11'b10110001001) ? 48'b101000110011000001000110000111010010111011010101 :
(key == 11'b10110001010) ? 48'b101000110010000110001010000111010000010001001001 :
(key == 11'b10110001011) ? 48'b101000110001001011010100000111001101100111010000 :
(key == 11'b10110001100) ? 48'b101000110000010000100001000111001010111101101011 :
(key == 11'b10110001101) ? 48'b101000101111010101110011000111001000010100011001 :
(key == 11'b10110001110) ? 48'b101000101110011011001000000111000101101011011011 :
(key == 11'b10110001111) ? 48'b101000101101100000100010000111000011000010110001 :
(key == 11'b10110010000) ? 48'b101000101100100110000000000111000000011010010111 :
(key == 11'b10110010001) ? 48'b101000101011101011100001000110111101110010010010 :
(key == 11'b10110010010) ? 48'b101000101010110001000110000110111011001010011110 :
(key == 11'b10110010011) ? 48'b101000101001110110110000000110111000100011000000 :
(key == 11'b10110010100) ? 48'b101000101000111100011101000110110101111011110001 :
(key == 11'b10110010101) ? 48'b101000101000000010001110000110110011010100110111 :
(key == 11'b10110010110) ? 48'b101000100111001000000011000110110000101110001111 :
(key == 11'b10110010111) ? 48'b101000100110001101111100000110101110000111111010 :
(key == 11'b10110011000) ? 48'b101000100101010011111000000110101011100001110110 :
(key == 11'b10110011001) ? 48'b101000100100011001111000000110101000111100000100 :
(key == 11'b10110011010) ? 48'b101000100011011111111110000110100110010110101001 :
(key == 11'b10110011011) ? 48'b101000100010100110000110000110100011110001011100 :
(key == 11'b10110011100) ? 48'b101000100001101100010010000110100001001100100011 :
(key == 11'b10110011101) ? 48'b101000100000110010100010000110011110100111111100 :
(key == 11'b10110011110) ? 48'b101000011111111000110110000110011100000011101010 :
(key == 11'b10110011111) ? 48'b101000011110111111001110000110011001011111100110 :
(key == 11'b10110100000) ? 48'b101000011110000101101010000110010110111011110111 :
(key == 11'b10110100001) ? 48'b101000011101001100001001000110010100011000011000 :
(key == 11'b10110100010) ? 48'b101000011100010010101100000110010001110101001101 :
(key == 11'b10110100011) ? 48'b101000011011011001010100000110001111010010010110 :
(key == 11'b10110100100) ? 48'b101000011010011111111111000110001100101111101100 :
(key == 11'b10110100101) ? 48'b101000011001100110101110000110001010001101010111 :
(key == 11'b10110100110) ? 48'b101000011000101101100000000110000111101011010011 :
(key == 11'b10110100111) ? 48'b101000010111110100010111000110000101001001100011 :
(key == 11'b10110101000) ? 48'b101000010110111011010001000110000010101000000011 :
(key == 11'b10110101001) ? 48'b101000010110000010010000000110000000000110110111 :
(key == 11'b10110101010) ? 48'b101000010101001001010000000101111101100101111000 :
(key == 11'b10110101011) ? 48'b101000010100010000010110000101111011000101001101 :
(key == 11'b10110101100) ? 48'b101000010011010111100000000101111000100100111000 :
(key == 11'b10110101101) ? 48'b101000010010011110101100000101110110000100101110 :
(key == 11'b10110101110) ? 48'b101000010001100101111100000101110011100100111000 :
(key == 11'b10110101111) ? 48'b101000010000101101010010000101110001000101010110 :
(key == 11'b10110110000) ? 48'b101000001111110100101010000101101110100110000010 :
(key == 11'b10110110001) ? 48'b101000001110111100000110000101101100000111000011 :
(key == 11'b10110110010) ? 48'b101000001110000011100110000101101001101000010011 :
(key == 11'b10110110011) ? 48'b101000001101001011001010000101100111001001110111 :
(key == 11'b10110110100) ? 48'b101000001100010010110000000101100100101011101000 :
(key == 11'b10110110101) ? 48'b101000001011011010011010000101100010001101101100 :
(key == 11'b10110110110) ? 48'b101000001010100010001001000101011111110000000010 :
(key == 11'b10110110111) ? 48'b101000001001101001111011000101011101010010101010 :
(key == 11'b10110111000) ? 48'b101000001000110001110001000101011010110101100010 :
(key == 11'b10110111001) ? 48'b101000000111111001101011000101011000011000101100 :
(key == 11'b10110111010) ? 48'b101000000111000001101000000101010101111100000111 :
(key == 11'b10110111011) ? 48'b101000000110001001101001000101010011011111110010 :
(key == 11'b10110111100) ? 48'b101000000101010001101110000101010001000011110000 :
(key == 11'b10110111101) ? 48'b101000000100011001110110000101001110100111111101 :
(key == 11'b10110111110) ? 48'b101000000011100010000010000101001100001100011011 :
(key == 11'b10110111111) ? 48'b101000000010101010010001000101001001110001001011 :
(key == 11'b10111000000) ? 48'b101000000001110010100100000101000111010110001011 :
(key == 11'b10111000001) ? 48'b101000000000111010111100000101000100111011011101 :
(key == 11'b10111000010) ? 48'b101000000000000011010110000101000010100000111110 :
(key == 11'b10111000011) ? 48'b100111111111001011110100000101000000000110110010 :
(key == 11'b10111000100) ? 48'b100111111110010100010110000100111101101100110110 :
(key == 11'b10111000101) ? 48'b100111111101011100111010000100111011010011001000 :
(key == 11'b10111000110) ? 48'b100111111100100101100011000100111000111001101101 :
(key == 11'b10111000111) ? 48'b100111111011101110010000000100110110100000100101 :
(key == 11'b10111001000) ? 48'b100111111010110111000000000100110100000111101000 :
(key == 11'b10111001001) ? 48'b100111111001111111110011000100110001101110111110 :
(key == 11'b10111001010) ? 48'b100111111001001000101011000100101111010110100111 :
(key == 11'b10111001011) ? 48'b100111111000010001100110000100101100111110011111 :
(key == 11'b10111001100) ? 48'b100111110111011010100100000100101010100110100110 :
(key == 11'b10111001101) ? 48'b100111110110100011100101000100101000001110111100 :
(key == 11'b10111001110) ? 48'b100111110101101100101010000100100101110111100101 :
(key == 11'b10111001111) ? 48'b100111110100110101110100000100100011100000100000 :
(key == 11'b10111010000) ? 48'b100111110011111111000001000100100001001001101001 :
(key == 11'b10111010001) ? 48'b100111110011001000010001000100011110110011000010 :
(key == 11'b10111010010) ? 48'b100111110010010001100100000100011100011100101100 :
(key == 11'b10111010011) ? 48'b100111110001011010111100000100011010000110100110 :
(key == 11'b10111010100) ? 48'b100111110000100100010110000100010111110000101101 :
(key == 11'b10111010101) ? 48'b100111101111101101110100000100010101011011000111 :
(key == 11'b10111010110) ? 48'b100111101110110111010110000100010011000101110010 :
(key == 11'b10111010111) ? 48'b100111101110000000111011000100010000110000101011 :
(key == 11'b10111011000) ? 48'b100111101101001010100011000100001110011011110011 :
(key == 11'b10111011001) ? 48'b100111101100010100010000000100001100000111001110 :
(key == 11'b10111011010) ? 48'b100111101011011101111111000100001001110010110111 :
(key == 11'b10111011011) ? 48'b100111101010100111110010000100000111011110110000 :
(key == 11'b10111011100) ? 48'b100111101001110001101000000100000101001010111000 :
(key == 11'b10111011101) ? 48'b100111101000111011100010000100000010110111010001 :
(key == 11'b10111011110) ? 48'b100111101000000101100000000100000000100011111000 :
(key == 11'b10111011111) ? 48'b100111100111001111100001000011111110010000110010 :
(key == 11'b10111100000) ? 48'b100111100110011001100101000011111011111101111000 :
(key == 11'b10111100001) ? 48'b100111100101100011101101000011111001101011010001 :
(key == 11'b10111100010) ? 48'b100111100100101101111000000011110111011000110110 :
(key == 11'b10111100011) ? 48'b100111100011111000000110000011110101000110101110 :
(key == 11'b10111100100) ? 48'b100111100011000010011000000011110010110100110011 :
(key == 11'b10111100101) ? 48'b100111100010001100101110000011110000100011001010 :
(key == 11'b10111100110) ? 48'b100111100001010111000111000011101110010001101110 :
(key == 11'b10111100111) ? 48'b100111100000100001100100000011101100000000100011 :
(key == 11'b10111101000) ? 48'b100111011111101100000011000011101001101111100110 :
(key == 11'b10111101001) ? 48'b100111011110110110100111000011100111011110111011 :
(key == 11'b10111101010) ? 48'b100111011110000001001100000011100101001110011011 :
(key == 11'b10111101011) ? 48'b100111011101001011110110000011100010111110001100 :
(key == 11'b10111101100) ? 48'b100111011100010110100100000011100000101110001100 :
(key == 11'b10111101101) ? 48'b100111011011100001010100000011011110011110011100 :
(key == 11'b10111101110) ? 48'b100111011010101100001000000011011100001110111011 :
(key == 11'b10111101111) ? 48'b100111011001110111000000000011011001111111101001 :
(key == 11'b10111110000) ? 48'b100111011001000001111010000011010111110000100110 :
(key == 11'b10111110001) ? 48'b100111011000001100111001000011010101100001110101 :
(key == 11'b10111110010) ? 48'b100111010111010111111010000011010011010011010000 :
(key == 11'b10111110011) ? 48'b100111010110100010111111000011010001000100111010 :
(key == 11'b10111110100) ? 48'b100111010101101110000111000011001110110110110011 :
(key == 11'b10111110101) ? 48'b100111010100111001010010000011001100101000111010 :
(key == 11'b10111110110) ? 48'b100111010100000100100001000011001010011011010001 :
(key == 11'b10111110111) ? 48'b100111010011001111110010000011001000001101110100 :
(key == 11'b10111111000) ? 48'b100111010010011011001000000011000110000000101001 :
(key == 11'b10111111001) ? 48'b100111010001100110100001000011000011110011101110 :
(key == 11'b10111111010) ? 48'b100111010000110001111101000011000001100111000001 :
(key == 11'b10111111011) ? 48'b100111001111111101011100000010111111011010100010 :
(key == 11'b10111111100) ? 48'b100111001111001000111110000010111101001110010000 :
(key == 11'b10111111101) ? 48'b100111001110010100100100000010111011000010001101 :
(key == 11'b10111111110) ? 48'b100111001101100000001101000010111000110110011001 :
(key == 11'b10111111111) ? 48'b100111001100101011111010000010110110101010110101 :
(key == 11'b11000000000) ? 48'b100111001011110111101001000010110100011111011111 :
(key == 11'b11000000001) ? 48'b100111001011000011011100000010110010010100010111 :
(key == 11'b11000000010) ? 48'b100111001010001111010010000010110000001001011111 :
(key == 11'b11000000011) ? 48'b100111001001011011001100000010101101111110110100 :
(key == 11'b11000000100) ? 48'b100111001000100111001000000010101011110100010111 :
(key == 11'b11000000101) ? 48'b100111000111110011001000000010101001101010001000 :
(key == 11'b11000000110) ? 48'b100111000110111111001011000010100111100000001000 :
(key == 11'b11000000111) ? 48'b100111000110001011010010000010100101010110010111 :
(key == 11'b11000001000) ? 48'b100111000101010111011100000010100011001100110100 :
(key == 11'b11000001001) ? 48'b100111000100100011101000000010100001000011100000 :
(key == 11'b11000001010) ? 48'b100111000011101111111000000010011110111010011001 :
(key == 11'b11000001011) ? 48'b100111000010111100001100000010011100110001100000 :
(key == 11'b11000001100) ? 48'b100111000010001000100010000010011010101000110100 :
(key == 11'b11000001101) ? 48'b100111000001010100111011000010011000100000011000 :
(key == 11'b11000001110) ? 48'b100111000000100001011000000010010110011000001010 :
(key == 11'b11000001111) ? 48'b100110111111101101111000000010010100010000001011 :
(key == 11'b11000010000) ? 48'b100110111110111010011100000010010010001000011001 :
(key == 11'b11000010001) ? 48'b100110111110000111000010000010010000000000110101 :
(key == 11'b11000010010) ? 48'b100110111101010011101100000010001101111001011111 :
(key == 11'b11000010011) ? 48'b100110111100100000011000000010001011110010010110 :
(key == 11'b11000010100) ? 48'b100110111011101101001000000010001001101011011010 :
(key == 11'b11000010101) ? 48'b100110111010111001111011000010000111100100101110 :
(key == 11'b11000010110) ? 48'b100110111010000110110010000010000101011110001111 :
(key == 11'b11000010111) ? 48'b100110111001010011101100000010000011011000000000 :
(key == 11'b11000011000) ? 48'b100110111000100000101000000010000001010001111100 :
(key == 11'b11000011001) ? 48'b100110110111101101100111000001111111001100000101 :
(key == 11'b11000011010) ? 48'b100110110110111010101010000001111101000110011110 :
(key == 11'b11000011011) ? 48'b100110110110000111110000000001111011000001000100 :
(key == 11'b11000011100) ? 48'b100110110101010100111001000001111000111011110111 :
(key == 11'b11000011101) ? 48'b100110110100100010000100000001110110110110110110 :
(key == 11'b11000011110) ? 48'b100110110011101111010100000001110100110010000110 :
(key == 11'b11000011111) ? 48'b100110110010111100100111000001110010101101100011 :
(key == 11'b11000100000) ? 48'b100110110010001001111100000001110000101001001110 :
(key == 11'b11000100001) ? 48'b100110110001010111010100000001101110100101000100 :
(key == 11'b11000100010) ? 48'b100110110000100100110000000001101100100001001000 :
(key == 11'b11000100011) ? 48'b100110101111110010001111000001101010011101011011 :
(key == 11'b11000100100) ? 48'b100110101110111111110001000001101000011001111010 :
(key == 11'b11000100101) ? 48'b100110101110001101010110000001100110010110100110 :
(key == 11'b11000100110) ? 48'b100110101101011010111110000001100100010011100010 :
(key == 11'b11000100111) ? 48'b100110101100101000101001000001100010010000101000 :
(key == 11'b11000101000) ? 48'b100110101011110110010110000001100000001101111100 :
(key == 11'b11000101001) ? 48'b100110101011000100001000000001011110001011011111 :
(key == 11'b11000101010) ? 48'b100110101010010001111100000001011100001001001111 :
(key == 11'b11000101011) ? 48'b100110101001011111110100000001011010000111001100 :
(key == 11'b11000101100) ? 48'b100110101000101101101110000001011000000101010100 :
(key == 11'b11000101101) ? 48'b100110100111111011101011000001010110000011101011 :
(key == 11'b11000101110) ? 48'b100110100111001001101100000001010100000010001111 :
(key == 11'b11000101111) ? 48'b100110100110010111110000000001010010000001000010 :
(key == 11'b11000110000) ? 48'b100110100101100101110110000001010000000000000000 :
(key == 11'b11000110001) ? 48'b100110100100110100000000000001001101111111001011 :
(key == 11'b11000110010) ? 48'b100110100100000010001100000001001011111110100001 :
(key == 11'b11000110011) ? 48'b100110100011010000011100000001001001111110001000 :
(key == 11'b11000110100) ? 48'b100110100010011110101110000001000111111101111010 :
(key == 11'b11000110101) ? 48'b100110100001101101000011000001000101111101110111 :
(key == 11'b11000110110) ? 48'b100110100000111011011100000001000011111110000100 :
(key == 11'b11000110111) ? 48'b100110100000001001111000000001000001111110011101 :
(key == 11'b11000111000) ? 48'b100110011111011000010110000000111111111111000010 :
(key == 11'b11000111001) ? 48'b100110011110100110111000000000111101111111110100 :
(key == 11'b11000111010) ? 48'b100110011101110101011100000000111100000000110011 :
(key == 11'b11000111011) ? 48'b100110011101000100000100000000111010000001111111 :
(key == 11'b11000111100) ? 48'b100110011100010010101110000000111000000011010110 :
(key == 11'b11000111101) ? 48'b100110011011100001011100000000110110000100111101 :
(key == 11'b11000111110) ? 48'b100110011010110000001100000000110100000110101111 :
(key == 11'b11000111111) ? 48'b100110011001111110111111000000110010001000101100 :
(key == 11'b11001000000) ? 48'b100110011001001101110110000000110000001010110111 :
(key == 11'b11001000001) ? 48'b100110011000011100101110000000101110001101001110 :
(key == 11'b11001000010) ? 48'b100110010111101011101010000000101100001111110001 :
(key == 11'b11001000011) ? 48'b100110010110111010101010000000101010010010100010 :
(key == 11'b11001000100) ? 48'b100110010110001001101100000000101000010101100000 :
(key == 11'b11001000101) ? 48'b100110010101011000110001000000100110011000101001 :
(key == 11'b11001000110) ? 48'b100110010100100111111001000000100100011011111111 :
(key == 11'b11001000111) ? 48'b100110010011110111000100000000100010011111100001 :
(key == 11'b11001001000) ? 48'b100110010011000110010000000000100000100011001110 :
(key == 11'b11001001001) ? 48'b100110010010010101100010000000011110100111001011 :
(key == 11'b11001001010) ? 48'b100110010001100100110101000000011100101011010001 :
(key == 11'b11001001011) ? 48'b100110010000110100001100000000011010101111101000 :
(key == 11'b11001001100) ? 48'b100110010000000011100110000000011000110100000111 :
(key == 11'b11001001101) ? 48'b100110001111010011000010000000010110111000110011 :
(key == 11'b11001001110) ? 48'b100110001110100010100000000000010100111101101011 :
(key == 11'b11001001111) ? 48'b100110001101110010000011000000010011000010110001 :
(key == 11'b11001010000) ? 48'b100110001101000001101000000000010001001000000000 :
(key == 11'b11001010001) ? 48'b100110001100010001010000000000001111001101011110 :
(key == 11'b11001010010) ? 48'b100110001011100000111010000000001101010011001000 :
(key == 11'b11001010011) ? 48'b100110001010110000101000000000001011011000111101 :
(key == 11'b11001010100) ? 48'b100110001010000000011000000000001001011110111101 :
(key == 11'b11001010101) ? 48'b100110001001010000001100000000000111100101001101 :
(key == 11'b11001010110) ? 48'b100110001000100000000010000000000101101011100101 :
(key == 11'b11001010111) ? 48'b100110000111101111111010000000000011110010001001 :
(key == 11'b11001011000) ? 48'b100110000110111111110110000000000001111000111011 :
(key == 11'b11001011001) ? 48'b100110000110001111110101011111111111111111110000 :
(key == 11'b11001011010) ? 48'b100110000101011111110110011111111100001110000011 :
(key == 11'b11001011011) ? 48'b100110000100101111111010011111111000011100101010 :
(key == 11'b11001011100) ? 48'b100110000100000000000010011111110100101011101110 :
(key == 11'b11001011101) ? 48'b100110000011010000001011011111110000111011000110 :
(key == 11'b11001011110) ? 48'b100110000010100000011000011111101101001010110111 :
(key == 11'b11001011111) ? 48'b100110000001110000100111011111101001011010111101 :
(key == 11'b11001100000) ? 48'b100110000001000000111001011111100101101011011011 :
(key == 11'b11001100001) ? 48'b100110000000010001001110011111100001111100010001 :
(key == 11'b11001100010) ? 48'b100101111111100001100110011111011110001101100000 :
(key == 11'b11001100011) ? 48'b100101111110110010000001011111011010011111000111 :
(key == 11'b11001100100) ? 48'b100101111110000010011111011111010110110001000111 :
(key == 11'b11001100101) ? 48'b100101111101010010111110011111010011000011011000 :
(key == 11'b11001100110) ? 48'b100101111100100011100010011111001111010110001000 :
(key == 11'b11001100111) ? 48'b100101111011110100001000011111001011101001001001 :
(key == 11'b11001101000) ? 48'b100101111011000100110000011111000111111100100010 :
(key == 11'b11001101001) ? 48'b100101111010010101011100011111000100010000010100 :
(key == 11'b11001101010) ? 48'b100101111001100110001010011111000000100100011101 :
(key == 11'b11001101011) ? 48'b100101111000110110111100011110111100111000111111 :
(key == 11'b11001101100) ? 48'b100101111000000111101111011110111001001101110010 :
(key == 11'b11001101101) ? 48'b100101110111011000100101011110110101100010111100 :
(key == 11'b11001101110) ? 48'b100101110110101001011110011110110001111000011111 :
(key == 11'b11001101111) ? 48'b100101110101111010011011011110101110001110011101 :
(key == 11'b11001110000) ? 48'b100101110101001011011010011110101010100100110000 :
(key == 11'b11001110001) ? 48'b100101110100011100011011011110100110111011010111 :
(key == 11'b11001110010) ? 48'b100101110011101101011110011110100011010010010010 :
(key == 11'b11001110011) ? 48'b100101110010111110100110011110011111101001101100 :
(key == 11'b11001110100) ? 48'b100101110010001111110000011110011100000001010111 :
(key == 11'b11001110101) ? 48'b100101110001100000111100011110011000011001010110 :
(key == 11'b11001110110) ? 48'b100101110000110010001010011110010100110001101101 :
(key == 11'b11001110111) ? 48'b100101110000000011011100011110010001001010011100 :
(key == 11'b11001111000) ? 48'b100101101111010100110001011110001101100011100010 :
(key == 11'b11001111001) ? 48'b100101101110100110001000011110001001111100111101 :
(key == 11'b11001111010) ? 48'b100101101101110111100010011110000110010110101111 :
(key == 11'b11001111011) ? 48'b100101101101001000111111011110000010110000111001 :
(key == 11'b11001111100) ? 48'b100101101100011010011110011101111111001011010011 :
(key == 11'b11001111101) ? 48'b100101101011101100000000011101111011100110001001 :
(key == 11'b11001111110) ? 48'b100101101010111101100101011101111000000001010110 :
(key == 11'b11001111111) ? 48'b100101101010001111001100011101110100011100110111 :
(key == 11'b11010000000) ? 48'b100101101001100000110110011101110000111000101000 :
(key == 11'b11010000001) ? 48'b100101101000110010100011011101101101010100111000 :
(key == 11'b11010000010) ? 48'b100101101000000100010010011101101001110001011001 :
(key == 11'b11010000011) ? 48'b100101100111010110000100011101100110001110010001 :
(key == 11'b11010000100) ? 48'b100101100110100111111001011101100010101011100000 :
(key == 11'b11010000101) ? 48'b100101100101111001110000011101011111001000111111 :
(key == 11'b11010000110) ? 48'b100101100101001011101010011101011011100110111001 :
(key == 11'b11010000111) ? 48'b100101100100011101100111011101011000000101001011 :
(key == 11'b11010001000) ? 48'b100101100011101111100110011101010100100011110000 :
(key == 11'b11010001001) ? 48'b100101100011000001101000011101010001000010100110 :
(key == 11'b11010001010) ? 48'b100101100010010011101100011101001101100001110010 :
(key == 11'b11010001011) ? 48'b100101100001100101110011011101001010000001011010 :
(key == 11'b11010001100) ? 48'b100101100000110111111101011101000110100001010101 :
(key == 11'b11010001101) ? 48'b100101100000001010001010011101000011000001100100 :
(key == 11'b11010001110) ? 48'b100101011111011100011010011100111111100010001101 :
(key == 11'b11010001111) ? 48'b100101011110101110101011011100111100000011000110 :
(key == 11'b11010010000) ? 48'b100101011110000000111110011100111000100100010000 :
(key == 11'b11010010001) ? 48'b100101011101010011010110011100110101000101110111 :
(key == 11'b11010010010) ? 48'b100101011100100101101111011100110001100111110010 :
(key == 11'b11010010011) ? 48'b100101011011111000001011011100101110001010000000 :
(key == 11'b11010010100) ? 48'b100101011011001010101010011100101010101100100010 :
(key == 11'b11010010101) ? 48'b100101011010011101001011011100100111001111011011 :
(key == 11'b11010010110) ? 48'b100101011001101111101111011100100011110010101011 :
(key == 11'b11010010111) ? 48'b100101011001000010010110011100100000010110001110 :
(key == 11'b11010011000) ? 48'b100101011000010100111110011100011100111010000000 :
(key == 11'b11010011001) ? 48'b100101010111100111101010011100011001011110010001 :
(key == 11'b11010011010) ? 48'b100101010110111010011001011100010110000010110101 :
(key == 11'b11010011011) ? 48'b100101010110001101001001011100010010100111101001 :
(key == 11'b11010011100) ? 48'b100101010101011111111101011100001111001100110111 :
(key == 11'b11010011101) ? 48'b100101010100110010110010011100001011110010010100 :
(key == 11'b11010011110) ? 48'b100101010100000101101011011100001000011000001001 :
(key == 11'b11010011111) ? 48'b100101010011011000100110011100000100111110010000 :
(key == 11'b11010100000) ? 48'b100101010010101011100011011100000001100100101011 :
(key == 11'b11010100001) ? 48'b100101010001111110100100011011111110001011100000 :
(key == 11'b11010100010) ? 48'b100101010001010001100110011011111010110010100100 :
(key == 11'b11010100011) ? 48'b100101010000100100101011011011110111011001111111 :
(key == 11'b11010100100) ? 48'b100101001111110111110010011011110100000001101101 :
(key == 11'b11010100101) ? 48'b100101001111001010111101011011110000101001110010 :
(key == 11'b11010100110) ? 48'b100101001110011110001010011011101101010010001001 :
(key == 11'b11010100111) ? 48'b100101001101110001011010011011101001111010110111 :
(key == 11'b11010101000) ? 48'b100101001101000100101100011011100110100011111000 :
(key == 11'b11010101001) ? 48'b100101001100010111111111011011100011001101001000 :
(key == 11'b11010101010) ? 48'b100101001011101011010110011011011111110110110010 :
(key == 11'b11010101011) ? 48'b100101001010111110101111011011011100100000101100 :
(key == 11'b11010101100) ? 48'b100101001010010010001100011011011001001010111111 :
(key == 11'b11010101101) ? 48'b100101001001100101101010011011010101110101100010 :
(key == 11'b11010101110) ? 48'b100101001000111001001010011011010010100000011011 :
(key == 11'b11010101111) ? 48'b100101001000001100101110011011001111001011101010 :
(key == 11'b11010110000) ? 48'b100101000111100000010100011011001011110111001001 :
(key == 11'b11010110001) ? 48'b100101000110110011111100011011001000100010111010 :
(key == 11'b11010110010) ? 48'b100101000110000111100110011011000101001111000001 :
(key == 11'b11010110011) ? 48'b100101000101011011010100011011000001111011011111 :
(key == 11'b11010110100) ? 48'b100101000100101111000100011010111110101000001100 :
(key == 11'b11010110101) ? 48'b100101000100000010110110011010111011010101010010 :
(key == 11'b11010110110) ? 48'b100101000011010110101011011010111000000010101000 :
(key == 11'b11010110111) ? 48'b100101000010101010100010011010110100110000010100 :
(key == 11'b11010111000) ? 48'b100101000001111110011100011010110001011110010010 :
(key == 11'b11010111001) ? 48'b100101000001010010011000011010101110001100100011 :
(key == 11'b11010111010) ? 48'b100101000000100110010110011010101010111011000110 :
(key == 11'b11010111011) ? 48'b100100111111111010010111011010100111101001111100 :
(key == 11'b11010111100) ? 48'b100100111111001110011011011010100100011001001011 :
(key == 11'b11010111101) ? 48'b100100111110100010100001011010100001001000101001 :
(key == 11'b11010111110) ? 48'b100100111101110110101001011010011101111000011010 :
(key == 11'b11010111111) ? 48'b100100111101001010110100011010011010101000100000 :
(key == 11'b11011000000) ? 48'b100100111100011111000010011010010111011000111100 :
(key == 11'b11011000001) ? 48'b100100111011110011010010011010010100001001101000 :
(key == 11'b11011000010) ? 48'b100100111011000111100010011010010000111010100010 :
(key == 11'b11011000011) ? 48'b100100111010011011110111011010001101101011110101 :
(key == 11'b11011000100) ? 48'b100100111001110000001110011010001010011101011011 :
(key == 11'b11011000101) ? 48'b100100111001000100101000011010000111001111010011 :
(key == 11'b11011000110) ? 48'b100100111000011001000100011010000100000001100000 :
(key == 11'b11011000111) ? 48'b100100110111101101100010011010000000110011111101 :
(key == 11'b11011001000) ? 48'b100100110111000010000010011001111101100110101111 :
(key == 11'b11011001001) ? 48'b100100110110010110100101011001111010011001110011 :
(key == 11'b11011001010) ? 48'b100100110101101011001010011001110111001101001010 :
(key == 11'b11011001011) ? 48'b100100110100111111110010011001110100000000110010 :
(key == 11'b11011001100) ? 48'b100100110100010100011100011001110000110100110000 :
(key == 11'b11011001101) ? 48'b100100110011101001001001011001101101101001000001 :
(key == 11'b11011001110) ? 48'b100100110010111101111000011001101010011101100011 :
(key == 11'b11011001111) ? 48'b100100110010010010101010011001100111010010011000 :
(key == 11'b11011010000) ? 48'b100100110001100111011110011001100100000111100010 :
(key == 11'b11011010001) ? 48'b100100110000111100010100011001100000111100111010 :
(key == 11'b11011010010) ? 48'b100100110000010001001100011001011101110010100101 :
(key == 11'b11011010011) ? 48'b100100101111100110000110011001011010101000100101 :
(key == 11'b11011010100) ? 48'b100100101110111011000100011001010111011110110110 :
(key == 11'b11011010101) ? 48'b100100101110010000000100011001010100010101011110 :
(key == 11'b11011010110) ? 48'b100100101101100101000110011001010001001100010100 :
(key == 11'b11011010111) ? 48'b100100101100111010001010011001001110000011011011 :
(key == 11'b11011011000) ? 48'b100100101100001111010000011001001010111010110100 :
(key == 11'b11011011001) ? 48'b100100101011100100011010011001000111110010100111 :
(key == 11'b11011011010) ? 48'b100100101010111001100110011001000100101010100111 :
(key == 11'b11011011011) ? 48'b100100101010001110110010011001000001100010110110 :
(key == 11'b11011011100) ? 48'b100100101001100100000010011000111110011011011010 :
(key == 11'b11011011101) ? 48'b100100101000111001010110011000111011010100010100 :
(key == 11'b11011011110) ? 48'b100100101000001110101010011000111000001101011011 :
(key == 11'b11011011111) ? 48'b100100100111100100000000011000110101000110110001 :
(key == 11'b11011100000) ? 48'b100100100110111001011010011000110010000000100000 :
(key == 11'b11011100001) ? 48'b100100100110001110110101011000101110111010011100 :
(key == 11'b11011100010) ? 48'b100100100101100100010011011000101011110100101110 :
(key == 11'b11011100011) ? 48'b100100100100111001110100011000101000101111010010 :
(key == 11'b11011100100) ? 48'b100100100100001111010110011000100101101010000111 :
(key == 11'b11011100101) ? 48'b100100100011100100111100011000100010100101001110 :
(key == 11'b11011100110) ? 48'b100100100010111010100010011000011111100000100010 :
(key == 11'b11011100111) ? 48'b100100100010010000001100011000011100011100010000 :
(key == 11'b11011101000) ? 48'b100100100001100101111000011000011001011000001011 :
(key == 11'b11011101001) ? 48'b100100100000111011100110011000010110010100011000 :
(key == 11'b11011101010) ? 48'b100100100000010001010110011000010011010000110110 :
(key == 11'b11011101011) ? 48'b100100011111100111001001011000010000001101100110 :
(key == 11'b11011101100) ? 48'b100100011110111100111110011000001101001010101000 :
(key == 11'b11011101101) ? 48'b100100011110010010110101011000001010000111111110 :
(key == 11'b11011101110) ? 48'b100100011101101000101110011000000111000101100010 :
(key == 11'b11011101111) ? 48'b100100011100111110101011011000000100000011011011 :
(key == 11'b11011110000) ? 48'b100100011100010100101000011000000001000001100010 :
(key == 11'b11011110001) ? 48'b100100011011101010101001010111111101111111111110 :
(key == 11'b11011110010) ? 48'b100100011011000000101100010111111010111110100111 :
(key == 11'b11011110011) ? 48'b100100011010010110110010010111110111111101101001 :
(key == 11'b11011110100) ? 48'b100100011001101100111000010111110100111100110101 :
(key == 11'b11011110101) ? 48'b100100011001000011000001010111110001111100010011 :
(key == 11'b11011110110) ? 48'b100100011000011001001100010111101110111100000010 :
(key == 11'b11011110111) ? 48'b100100010111101111011100010111101011111100001000 :
(key == 11'b11011111000) ? 48'b100100010111000101101011010111101000111100011010 :
(key == 11'b11011111001) ? 48'b100100010110011011111101010111100101111100111100 :
(key == 11'b11011111010) ? 48'b100100010101110010010010010111100010111101110000 :
(key == 11'b11011111011) ? 48'b100100010101001000101010010111011111111110111011 :
(key == 11'b11011111100) ? 48'b100100010100011111000010010111011101000000010001 :
(key == 11'b11011111101) ? 48'b100100010011110101011101010111011010000001111000 :
(key == 11'b11011111110) ? 48'b100100010011001011111010010111010111000011110000 :
(key == 11'b11011111111) ? 48'b100100010010100010011100010111010100000110000000 :
(key == 11'b11100000000) ? 48'b100100010001111000111101010111010001001000011011 :
(key == 11'b11100000001) ? 48'b100100010001001111100001010111001110001011000110 :
(key == 11'b11100000010) ? 48'b100100010000100110001000010111001011001110000010 :
(key == 11'b11100000011) ? 48'b100100001111111100110000010111001000010001010000 :
(key == 11'b11100000100) ? 48'b100100001111010011011100010111000101010100110010 :
(key == 11'b11100000101) ? 48'b100100001110101010001000010111000010011000100001 :
(key == 11'b11100000110) ? 48'b100100001110000000111000010110111111011100100001 :
(key == 11'b11100000111) ? 48'b100100001101010111101001010110111100100000110010 :
(key == 11'b11100001000) ? 48'b100100001100101110011101010110111001100101010100 :
(key == 11'b11100001001) ? 48'b100100001100000101010011010110110110101010001000 :
(key == 11'b11100001010) ? 48'b100100001011011100001011010110110011101111001100 :
(key == 11'b11100001011) ? 48'b100100001010110011000101010110110000110100011101 :
(key == 11'b11100001100) ? 48'b100100001010001010000010010110101101111010000010 :
(key == 11'b11100001101) ? 48'b100100001001100001000000010110101010111111110110 :
(key == 11'b11100001110) ? 48'b100100001000111000000001010110101000000101111100 :
(key == 11'b11100001111) ? 48'b100100001000001111000100010110100101001100010001 :
(key == 11'b11100010000) ? 48'b100100000111100110001001010110100010010010110110 :
(key == 11'b11100010001) ? 48'b100100000110111101010001010110011111011001110000 :
(key == 11'b11100010010) ? 48'b100100000110010100011010010110011100100000110111 :
(key == 11'b11100010011) ? 48'b100100000101101011100110010110011001101000001011 :
(key == 11'b11100010100) ? 48'b100100000101000010110100010110010110101111110100 :
(key == 11'b11100010101) ? 48'b100100000100011010000100010110010011110111101100 :
(key == 11'b11100010110) ? 48'b100100000011110001010110010110010000111111110011 :
(key == 11'b11100010111) ? 48'b100100000011001000101010010110001110001000001101 :
(key == 11'b11100011000) ? 48'b100100000010100000000000010110001011010000110100 :
(key == 11'b11100011001) ? 48'b100100000001110111011001010110001000011001101100 :
(key == 11'b11100011010) ? 48'b100100000001001110110100010110000101100010111000 :
(key == 11'b11100011011) ? 48'b100100000000100110010010010110000010101100010010 :
(key == 11'b11100011100) ? 48'b100011111111111101110001010101111111110101111100 :
(key == 11'b11100011101) ? 48'b100011111111010101010010010101111100111111110010 :
(key == 11'b11100011110) ? 48'b100011111110101100110100010101111010001001111010 :
(key == 11'b11100011111) ? 48'b100011111110000100011010010101110111010100010101 :
(key == 11'b11100100000) ? 48'b100011111101011100000010010101110100011110111110 :
(key == 11'b11100100001) ? 48'b100011111100110011101011010101110001101001110011 :
(key == 11'b11100100010) ? 48'b100011111100001011010111010101101110110100111100 :
(key == 11'b11100100011) ? 48'b100011111011100011000101010101101100000000010110 :
(key == 11'b11100100100) ? 48'b100011111010111010110101010101101001001011111101 :
(key == 11'b11100100101) ? 48'b100011111010010010100111010101100110010111110100 :
(key == 11'b11100100110) ? 48'b100011111001101010011100010101100011100011111111 :
(key == 11'b11100100111) ? 48'b100011111001000010010010010101100000110000010111 :
(key == 11'b11100101000) ? 48'b100011111000011010001010010101011101111100111100 :
(key == 11'b11100101001) ? 48'b100011110111110010000110010101011011001001110100 :
(key == 11'b11100101010) ? 48'b100011110111001010000010010101011000010110111010 :
(key == 11'b11100101011) ? 48'b100011110110100010000001010101010101100100010000 :
(key == 11'b11100101100) ? 48'b100011110101111010000010010101010010110001110110 :
(key == 11'b11100101101) ? 48'b100011110101010010000101010101001111111111101100 :
(key == 11'b11100101110) ? 48'b100011110100101010001001010101001101001101101100 :
(key == 11'b11100101111) ? 48'b100011110100000010010001010101001010011100000010 :
(key == 11'b11100110000) ? 48'b100011110011011010011010010101000111101010100110 :
(key == 11'b11100110001) ? 48'b100011110010110010100110010101000100111001011010 :
(key == 11'b11100110010) ? 48'b100011110010001010110010010101000010001000011011 :
(key == 11'b11100110011) ? 48'b100011110001100011000010010100111111010111101011 :
(key == 11'b11100110100) ? 48'b100011110000111011010011010100111100100111001100 :
(key == 11'b11100110101) ? 48'b100011110000010011100111010100111001110110111110 :
(key == 11'b11100110110) ? 48'b100011101111101011111101010100110111000110111110 :
(key == 11'b11100110111) ? 48'b100011101111000100010100010100110100010111001100 :
(key == 11'b11100111000) ? 48'b100011101110011100101110010100110001100111101010 :
(key == 11'b11100111001) ? 48'b100011101101110101001010010100101110111000010101 :
(key == 11'b11100111010) ? 48'b100011101101001101101000010100101100001001010011 :
(key == 11'b11100111011) ? 48'b100011101100100110001000010100101001011010011110 :
(key == 11'b11100111100) ? 48'b100011101011111110101010010100100110101011111000 :
(key == 11'b11100111101) ? 48'b100011101011010111001110010100100011111101100011 :
(key == 11'b11100111110) ? 48'b100011101010101111110100010100100001001111011010 :
(key == 11'b11100111111) ? 48'b100011101010001000011100010100011110100001100010 :
(key == 11'b11101000000) ? 48'b100011101001100001000110010100011011110011111100 :
(key == 11'b11101000001) ? 48'b100011101000111001110011010100011001000110100011 :
(key == 11'b11101000010) ? 48'b100011101000010010100001010100010110011001010110 :
(key == 11'b11101000011) ? 48'b100011100111101011010000010100010011101100010111 :
(key == 11'b11101000100) ? 48'b100011100111000100000011010100010000111111101010 :
(key == 11'b11101000101) ? 48'b100011100110011100110111010100001110010011001010 :
(key == 11'b11101000110) ? 48'b100011100101110101101101010100001011100110111010 :
(key == 11'b11101000111) ? 48'b100011100101001110100110010100001000111010111010 :
(key == 11'b11101001000) ? 48'b100011100100100111100000010100000110001111001001 :
(key == 11'b11101001001) ? 48'b100011100100000000011100010100000011100011100010 :
(key == 11'b11101001010) ? 48'b100011100011011001011010010100000000111000001101 :
(key == 11'b11101001011) ? 48'b100011100010110010011010010011111110001101000101 :
(key == 11'b11101001100) ? 48'b100011100010001011011110010011111011100010010000 :
(key == 11'b11101001101) ? 48'b100011100001100100100010010011111000110111101000 :
(key == 11'b11101001110) ? 48'b100011100000111101101000010011110110001101001100 :
(key == 11'b11101001111) ? 48'b100011100000010110110000010011110011100011000000 :
(key == 11'b11101010000) ? 48'b100011011111101111111010010011110000111001000000 :
(key == 11'b11101010001) ? 48'b100011011111001001000111010011101110001111010010 :
(key == 11'b11101010010) ? 48'b100011011110100010010101010011101011100101110010 :
(key == 11'b11101010011) ? 48'b100011011101111011100110010011101000111100100000 :
(key == 11'b11101010100) ? 48'b100011011101010100111000010011100110010011011100 :
(key == 11'b11101010101) ? 48'b100011011100101110001100010011100011101010101010 :
(key == 11'b11101010110) ? 48'b100011011100000111100010010011100001000010000001 :
(key == 11'b11101010111) ? 48'b100011011011100000111010010011011110011001101000 :
(key == 11'b11101011000) ? 48'b100011011010111010010100010011011011110001011110 :
(key == 11'b11101011001) ? 48'b100011011010010011110001010011011001001001100100 :
(key == 11'b11101011010) ? 48'b100011011001101101001111010011010110100001110110 :
(key == 11'b11101011011) ? 48'b100011011001000110101111010011010011111010010111 :
(key == 11'b11101011100) ? 48'b100011011000100000010001010011010001010011000101 :
(key == 11'b11101011101) ? 48'b100011010111111001110101010011001110101100000010 :
(key == 11'b11101011110) ? 48'b100011010111010011011011010011001100000101001110 :
(key == 11'b11101011111) ? 48'b100011010110101101000011010011001001011110100111 :
(key == 11'b11101100000) ? 48'b100011010110000110101101010011000110111000001111 :
(key == 11'b11101100001) ? 48'b100011010101100000011001010011000100010010000110 :
(key == 11'b11101100010) ? 48'b100011010100111010000111010011000001101100001010 :
(key == 11'b11101100011) ? 48'b100011010100010011110110010010111111000110010111 :
(key == 11'b11101100100) ? 48'b100011010011101101101000010010111100100000111001 :
(key == 11'b11101100101) ? 48'b100011010011000111011100010010111001111011101000 :
(key == 11'b11101100110) ? 48'b100011010010100001010010010010110111010110100110 :
(key == 11'b11101100111) ? 48'b100011010001111011001001010010110100110001101111 :
(key == 11'b11101101000) ? 48'b100011010001010101000010010010110010001101000101 :
(key == 11'b11101101001) ? 48'b100011010000101110111110010010101111101000101110 :
(key == 11'b11101101010) ? 48'b100011010000001000111011010010101101000100011110 :
(key == 11'b11101101011) ? 48'b100011001111100010111001010010101010100000011100 :
(key == 11'b11101101100) ? 48'b100011001110111100111010010010100111111100101100 :
(key == 11'b11101101101) ? 48'b100011001110010110111110010010100101011001001010 :
(key == 11'b11101101110) ? 48'b100011001101110001000100010010100010110101111000 :
(key == 11'b11101101111) ? 48'b100011001101001011001010010010100000010010101111 :
(key == 11'b11101110000) ? 48'b100011001100100101010010010010011101101111110010 :
(key == 11'b11101110001) ? 48'b100011001011111111011101010010011011001101000111 :
(key == 11'b11101110010) ? 48'b100011001011011001101010010010011000101010101000 :
(key == 11'b11101110011) ? 48'b100011001010110011111000010010010110001000010100 :
(key == 11'b11101110100) ? 48'b100011001010001110001000010010010011100110010100 :
(key == 11'b11101110101) ? 48'b100011001001101000011010010010010001000100011100 :
(key == 11'b11101110110) ? 48'b100011001001000010101110010010001110100010110010 :
(key == 11'b11101110111) ? 48'b100011001000011101000100010010001100000001011000 :
(key == 11'b11101111000) ? 48'b100011000111110111011101010010001001100000001110 :
(key == 11'b11101111001) ? 48'b100011000111010001110110010010000110111111001011 :
(key == 11'b11101111010) ? 48'b100011000110101100010010010010000100011110011000 :
(key == 11'b11101111011) ? 48'b100011000110000110110000010010000001111101110100 :
(key == 11'b11101111100) ? 48'b100011000101100001010000010001111111011101011110 :
(key == 11'b11101111101) ? 48'b100011000100111011110001010001111100111101010100 :
(key == 11'b11101111110) ? 48'b100011000100010110010100010001111010011101010111 :
(key == 11'b11101111111) ? 48'b100011000011110000111000010001110111111101100100 :
(key == 11'b11110000000) ? 48'b100011000011001011100000010001110101011110000100 :
(key == 11'b11110000001) ? 48'b100011000010100110001000010001110010111110101101 :
(key == 11'b11110000010) ? 48'b100011000010000000110011010001110000011111100100 :
(key == 11'b11110000011) ? 48'b100011000001011011100000010001101110000000101011 :
(key == 11'b11110000100) ? 48'b100011000000110110001110010001101011100010000000 :
(key == 11'b11110000101) ? 48'b100011000000010000111111010001101001000011100001 :
(key == 11'b11110000110) ? 48'b100010111111101011110001010001100110100101001101 :
(key == 11'b11110000111) ? 48'b100010111111000110100100010001100100000111000101 :
(key == 11'b11110001000) ? 48'b100010111110100001011010010001100001101001001100 :
(key == 11'b11110001001) ? 48'b100010111101111100010010010001011111001011011110 :
(key == 11'b11110001010) ? 48'b100010111101010111001011010001011100101110000000 :
(key == 11'b11110001011) ? 48'b100010111100110010000111010001011010010000110000 :
(key == 11'b11110001100) ? 48'b100010111100001101000100010001010111110011101100 :
(key == 11'b11110001101) ? 48'b100010111011101000000100010001010101010110110110 :
(key == 11'b11110001110) ? 48'b100010111011000011000100010001010010111010001100 :
(key == 11'b11110001111) ? 48'b100010111010011110000111010001010000011101101101 :
(key == 11'b11110010000) ? 48'b100010111001111001001011010001001110000001011010 :
(key == 11'b11110010001) ? 48'b100010111001010100010010010001001011100101011001 :
(key == 11'b11110010010) ? 48'b100010111000101111011010010001001001001001100100 :
(key == 11'b11110010011) ? 48'b100010111000001010100100010001000110101101111001 :
(key == 11'b11110010100) ? 48'b100010110111100101110000010001000100010010011011 :
(key == 11'b11110010101) ? 48'b100010110111000000111110010001000001110111001010 :
(key == 11'b11110010110) ? 48'b100010110110011100001101010000111111011100000110 :
(key == 11'b11110010111) ? 48'b100010110101110111011110010000111101000001010000 :
(key == 11'b11110011000) ? 48'b100010110101010010110010010000111010100110100101 :
(key == 11'b11110011001) ? 48'b100010110100101110000110010000111000001100000110 :
(key == 11'b11110011010) ? 48'b100010110100001001011110010000110101110001111000 :
(key == 11'b11110011011) ? 48'b100010110011100100110110010000110011010111110011 :
(key == 11'b11110011100) ? 48'b100010110011000000010000010000110000111101111100 :
(key == 11'b11110011101) ? 48'b100010110010011011101101010000101110100100010100 :
(key == 11'b11110011110) ? 48'b100010110001110111001010010000101100001010110100 :
(key == 11'b11110011111) ? 48'b100010110001010010101011010000101001110001100101 :
(key == 11'b11110100000) ? 48'b100010110000101110001100010000100111011000011111 :
(key == 11'b11110100001) ? 48'b100010110000001001101111010000100100111111100100 :
(key == 11'b11110100010) ? 48'b100010101111100101010100010000100010100110110111 :
(key == 11'b11110100011) ? 48'b100010101111000000111011010000100000001110011001 :
(key == 11'b11110100100) ? 48'b100010101110011100100100010000011101110110000110 :
(key == 11'b11110100101) ? 48'b100010101101111000001110010000011011011101111110 :
(key == 11'b11110100110) ? 48'b100010101101010011111010010000011001000110000010 :
(key == 11'b11110100111) ? 48'b100010101100101111101000010000010110101110010100 :
(key == 11'b11110101000) ? 48'b100010101100001011011000010000010100010110110101 :
(key == 11'b11110101001) ? 48'b100010101011100111001010010000010001111111100000 :
(key == 11'b11110101010) ? 48'b100010101011000010111110010000001111101000011010 :
(key == 11'b11110101011) ? 48'b100010101010011110110100010000001101010001011111 :
(key == 11'b11110101100) ? 48'b100010101001111010101010010000001010111010110000 :
(key == 11'b11110101101) ? 48'b100010101001010110100011010000001000100100001011 :
(key == 11'b11110101110) ? 48'b100010101000110010011101010000000110001101110010 :
(key == 11'b11110101111) ? 48'b100010101000001110011001010000000011110111100111 :
(key == 11'b11110110000) ? 48'b100010100111101010010111010000000001100001100111 :
(key == 11'b11110110001) ? 48'b100010100111000110010111001111111111001011110101 :
(key == 11'b11110110010) ? 48'b100010100110100010011000001111111100110110001110 :
(key == 11'b11110110011) ? 48'b100010100101111110011100001111111010100000110010 :
(key == 11'b11110110100) ? 48'b100010100101011010100001001111111000001011100101 :
(key == 11'b11110110101) ? 48'b100010100100110110101000001111110101110110100011 :
(key == 11'b11110110110) ? 48'b100010100100010010110000001111110011100001101111 :
(key == 11'b11110110111) ? 48'b100010100011101110111010001111110001001101000010 :
(key == 11'b11110111000) ? 48'b100010100011001011000110001111101110111000100100 :
(key == 11'b11110111001) ? 48'b100010100010100111010100001111101100100100010101 :
(key == 11'b11110111010) ? 48'b100010100010000011100100001111101010010000001101 :
(key == 11'b11110111011) ? 48'b100010100001011111110100001111100111111100010000 :
(key == 11'b11110111100) ? 48'b100010100000111100001000001111100101101000100100 :
(key == 11'b11110111101) ? 48'b100010100000011000011100001111100011010101000011 :
(key == 11'b11110111110) ? 48'b100010011111110100110011001111100001000001101101 :
(key == 11'b11110111111) ? 48'b100010011111010001001011001111011110101110100010 :
(key == 11'b11111000000) ? 48'b100010011110101101100100001111011100011011100010 :
(key == 11'b11111000001) ? 48'b100010011110001010000000001111011010001000101101 :
(key == 11'b11111000010) ? 48'b100010011101100110011101001111010111110110000110 :
(key == 11'b11111000011) ? 48'b100010011101000010111100001111010101100011101010 :
(key == 11'b11111000100) ? 48'b100010011100011111011100001111010011010001011100 :
(key == 11'b11111000101) ? 48'b100010011011111011111111001111010000111111011000 :
(key == 11'b11111000110) ? 48'b100010011011011000100011001111001110101101100000 :
(key == 11'b11111000111) ? 48'b100010011010110101001000001111001100011011110010 :
(key == 11'b11111001000) ? 48'b100010011010010001110000001111001010001010010011 :
(key == 11'b11111001001) ? 48'b100010011001101110011010001111000111111000111110 :
(key == 11'b11111001010) ? 48'b100010011001001011000100001111000101100111110100 :
(key == 11'b11111001011) ? 48'b100010011000100111110000001111000011010110110101 :
(key == 11'b11111001100) ? 48'b100010011000000100011111001111000001000110000100 :
(key == 11'b11111001101) ? 48'b100010010111100001001111001110111110110101011101 :
(key == 11'b11111001110) ? 48'b100010010110111110000001001110111100100101000100 :
(key == 11'b11111001111) ? 48'b100010010110011010110101001110111010010100110110 :
(key == 11'b11111010000) ? 48'b100010010101110111101010001110111000000100110000 :
(key == 11'b11111010001) ? 48'b100010010101010100100001001110110101110100111100 :
(key == 11'b11111010010) ? 48'b100010010100110001011001001110110011100101001110 :
(key == 11'b11111010011) ? 48'b100010010100001110010011001110110001010101101011 :
(key == 11'b11111010100) ? 48'b100010010011101011001111001110101111000110010110 :
(key == 11'b11111010101) ? 48'b100010010011001000001100001110101100110111001100 :
(key == 11'b11111010110) ? 48'b100010010010100101001100001110101010101000001100 :
(key == 11'b11111010111) ? 48'b100010010010000010001100001110101000011001010110 :
(key == 11'b11111011000) ? 48'b100010010001011111010000001110100110001010110010 :
(key == 11'b11111011001) ? 48'b100010010000111100010100001110100011111100010110 :
(key == 11'b11111011010) ? 48'b100010010000011001011010001110100001101110000100 :
(key == 11'b11111011011) ? 48'b100010001111110110100001001110011111011111111100 :
(key == 11'b11111011100) ? 48'b100010001111010011101010001110011101010010000000 :
(key == 11'b11111011101) ? 48'b100010001110110000110100001110011011000100010001 :
(key == 11'b11111011110) ? 48'b100010001110001110000001001110011000110110101100 :
(key == 11'b11111011111) ? 48'b100010001101101011010000001110010110101001010110 :
(key == 11'b11111100000) ? 48'b100010001101001000100000001110010100011100001010 :
(key == 11'b11111100001) ? 48'b100010001100100101110001001110010010001111000101 :
(key == 11'b11111100010) ? 48'b100010001100000011000100001110010000000010001110 :
(key == 11'b11111100011) ? 48'b100010001011100000011001001110001101110101100010 :
(key == 11'b11111100100) ? 48'b100010001010111101110000001110001011101001000010 :
(key == 11'b11111100101) ? 48'b100010001010011011001000001110001001011100101011 :
(key == 11'b11111100110) ? 48'b100010001001111000100001001110000111010000011110 :
(key == 11'b11111100111) ? 48'b100010001001010101111100001110000101000100011111 :
(key == 11'b11111101000) ? 48'b100010001000110011011010001110000010111000101010 :
(key == 11'b11111101001) ? 48'b100010001000010000111000001110000000101101000000 :
(key == 11'b11111101010) ? 48'b100010000111101110011000001101111110100001100000 :
(key == 11'b11111101011) ? 48'b100010000111001011111010001101111100010110001101 :
(key == 11'b11111101100) ? 48'b100010000110101001011110001101111010001011000101 :
(key == 11'b11111101101) ? 48'b100010000110000111000011001101111000000000001000 :
(key == 11'b11111101110) ? 48'b100010000101100100101010001101110101110101010100 :
(key == 11'b11111101111) ? 48'b100010000101000010010011001101110011101010101111 :
(key == 11'b11111110000) ? 48'b100010000100011111111101001101110001100000010001 :
(key == 11'b11111110001) ? 48'b100010000011111101101000001101101111010101111101 :
(key == 11'b11111110010) ? 48'b100010000011011011010110001101101101001011110110 :
(key == 11'b11111110011) ? 48'b100010000010111001000100001101101011000001111010 :
(key == 11'b11111110100) ? 48'b100010000010010110110101001101101000111000001000 :
(key == 11'b11111110101) ? 48'b100010000001110100100111001101100110101110100010 :
(key == 11'b11111110110) ? 48'b100010000001010010011010001101100100100101000100 :
(key == 11'b11111110111) ? 48'b100010000000110000010000001101100010011011110101 :
(key == 11'b11111111000) ? 48'b100010000000001110001000001101100000010010110000 :
(key == 11'b11111111001) ? 48'b100001111111101100000000001101011110001001110010 :
(key == 11'b11111111010) ? 48'b100001111111001001111010001101011100000001000001 :
(key == 11'b11111111011) ? 48'b100001111110100111110110001101011001111000011010 :
(key == 11'b11111111100) ? 48'b100001111110000101110100001101010111110000000010 :
(key == 11'b11111111101) ? 48'b100001111101100011110010001101010101100111110000 :
(key == 11'b11111111110) ? 48'b100001111101000001110010001101010011011111101000 :
(key == 11'b11111111111) ? 48'b100001111100011111110101001101010001010111101110 : 48'd0;

endmodule

`default_nettype wire
