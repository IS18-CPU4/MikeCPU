`default_nettype none

module fsqrt
   ( input wire [31:0] x,
     output wire [31:0] y,
     output wire ovf);

   // split sequence to each subsequence
   wire xs;
   wire [7:0] xe;
   wire [22:0] xm;
   assign {xs, xe, xm} = x;

   // calc s
   wire s;
   assign s = xs;

   wire [7:0] shift_xe;
   assign shift_xe = xe >> 1;

   // calc e
   wire [7:0] e;
   assign e = (xe[0] == 1) ? 8'd189 - shift_xe : 8'd190 - shift_xe; 

   // calc m
   wire [22:0] m;
   wire [45:0] val;
   wire [10:0] key;
   assign key = {xe[0], xm[22:13]};
   // lookup table and get constant and grad
   lookup_table lt(key, val);
   wire [22:0] constant;
   wire [22:0] grad;
   // constant supplements 1 at the MSB
   assign constant = val[45:23];
   assign grad = val[22:0];
   wire [45:0] grad2;
   assign grad2 = xm * grad;
   assign m = constant - grad2;

   wire [31:0] tmp_y;
   fmul u1(x, {s, e, m}, tmp_y, ovf);

   wire [31:0] root2;
   assign root2 = 31'b00111111101101010000010011110011;

   wire [7:0] odd_zero_ye;
   assign odd_zero_ye = shift_xe + 8'd64;

   wire [31:0] even_zero_y;
   wire [7:0] even_zero_tmp_ye;
   assign even_zero_y = 8'd63 + shift_xe;
   wire tmp_ovf;
   fmul u2(root2, {xs, even_zero_tmp_ye, xm}, even_zero_y, tmp_ovf);

   assign y = (xm != 23'd0) ? tmp_y :
              (xe[0] == 1) ? {xs, odd_zero_ye, xm} : even_zero_y;

endmodule

module lookup_table
   ( input wire [10:0] key,
     output wire [45:0] value);

   assign value =
(key == 11'b00000000000) ? 46'b0000111101110110011110000001111011101100111100 :
(key == 11'b00000000001) ? 46'b0000111101010100100101000001111010101001001010 :
(key == 11'b00000000010) ? 46'b0000111100110010101111000001111001100101011110 :
(key == 11'b00000000011) ? 46'b0000111100010000111100000001111000100001111000 :
(key == 11'b00000000100) ? 46'b0000111011101111001100100001110111011110011001 :
(key == 11'b00000000101) ? 46'b0000111011001101100000000001110110011011000000 :
(key == 11'b00000000110) ? 46'b0000111010101011110111000001110101010111101110 :
(key == 11'b00000000111) ? 46'b0000111010001010010001000001110100010100100010 :
(key == 11'b00000001000) ? 46'b0000111001101000101101100001110011010001011011 :
(key == 11'b00000001001) ? 46'b0000111001000111001110000001110010001110011100 :
(key == 11'b00000001010) ? 46'b0000111000100101110001000001110001001011100010 :
(key == 11'b00000001011) ? 46'b0000111000000100010111100001110000001000101111 :
(key == 11'b00000001100) ? 46'b0000110111100011000001000001101111000110000010 :
(key == 11'b00000001101) ? 46'b0000110111000001101101100001101110000011011011 :
(key == 11'b00000001110) ? 46'b0000110110100000011101000001101101000000111010 :
(key == 11'b00000001111) ? 46'b0000110101111111001111100001101011111110011111 :
(key == 11'b00000010000) ? 46'b0000110101011110000101000001101010111100001010 :
(key == 11'b00000010001) ? 46'b0000110100111100111110000001101001111001111100 :
(key == 11'b00000010010) ? 46'b0000110100011011111010000001101000110111110100 :
(key == 11'b00000010011) ? 46'b0000110011111010111001000001100111110101110010 :
(key == 11'b00000010100) ? 46'b0000110011011001111011000001100110110011110110 :
(key == 11'b00000010101) ? 46'b0000110010111000111111100001100101110001111111 :
(key == 11'b00000010110) ? 46'b0000110010011000000111000001100100110000001110 :
(key == 11'b00000010111) ? 46'b0000110001110111010010000001100011101110100100 :
(key == 11'b00000011000) ? 46'b0000110001010110100000000001100010101101000000 :
(key == 11'b00000011001) ? 46'b0000110000110101110001000001100001101011100010 :
(key == 11'b00000011010) ? 46'b0000110000010101000101100001100000101010001011 :
(key == 11'b00000011011) ? 46'b0000101111110100011100000001011111101000111000 :
(key == 11'b00000011100) ? 46'b0000101111010011110110000001011110100111101100 :
(key == 11'b00000011101) ? 46'b0000101110110011010010100001011101100110100101 :
(key == 11'b00000011110) ? 46'b0000101110010010110011000001011100100101100110 :
(key == 11'b00000011111) ? 46'b0000101101110010010101100001011011100100101011 :
(key == 11'b00000100000) ? 46'b0000101101010001111011000001011010100011110110 :
(key == 11'b00000100001) ? 46'b0000101100110001100100000001011001100011001000 :
(key == 11'b00000100010) ? 46'b0000101100010001001111100001011000100010011111 :
(key == 11'b00000100011) ? 46'b0000101011110000111110100001010111100001111101 :
(key == 11'b00000100100) ? 46'b0000101011010000110000000001010110100001100000 :
(key == 11'b00000100101) ? 46'b0000101010110000100100000001010101100001001000 :
(key == 11'b00000100110) ? 46'b0000101010010000011011100001010100100000110111 :
(key == 11'b00000100111) ? 46'b0000101001110000010110000001010011100000101100 :
(key == 11'b00000101000) ? 46'b0000101001010000010010100001010010100000100101 :
(key == 11'b00000101001) ? 46'b0000101000110000010010100001010001100000100101 :
(key == 11'b00000101010) ? 46'b0000101000010000010101100001010000100000101011 :
(key == 11'b00000101011) ? 46'b0000100111110000011011000001001111100000110110 :
(key == 11'b00000101100) ? 46'b0000100111010000100100000001001110100001001000 :
(key == 11'b00000101101) ? 46'b0000100110110000101111000001001101100001011110 :
(key == 11'b00000101110) ? 46'b0000100110010000111101100001001100100001111011 :
(key == 11'b00000101111) ? 46'b0000100101110001001111000001001011100010011110 :
(key == 11'b00000110000) ? 46'b0000100101010001100011000001001010100011000110 :
(key == 11'b00000110001) ? 46'b0000100100110001111001100001001001100011110011 :
(key == 11'b00000110010) ? 46'b0000100100010010010011000001001000100100100110 :
(key == 11'b00000110011) ? 46'b0000100011110010110000000001000111100101100000 :
(key == 11'b00000110100) ? 46'b0000100011010011001111000001000110100110011110 :
(key == 11'b00000110101) ? 46'b0000100010110011110001100001000101100111100011 :
(key == 11'b00000110110) ? 46'b0000100010010100010110000001000100101000101100 :
(key == 11'b00000110111) ? 46'b0000100001110100111110000001000011101001111100 :
(key == 11'b00000111000) ? 46'b0000100001010101101000000001000010101011010000 :
(key == 11'b00000111001) ? 46'b0000100000110110010110000001000001101100101100 :
(key == 11'b00000111010) ? 46'b0000100000010111000110000001000000101110001100 :
(key == 11'b00000111011) ? 46'b0000011111110111111000100000111111101111110001 :
(key == 11'b00000111100) ? 46'b0000011111011000101110000000111110110001011100 :
(key == 11'b00000111101) ? 46'b0000011110111001100111000000111101110011001110 :
(key == 11'b00000111110) ? 46'b0000011110011010100010000000111100110101000100 :
(key == 11'b00000111111) ? 46'b0000011101111011100000000000111011110111000000 :
(key == 11'b00001000000) ? 46'b0000011101011100100000100000111010111001000001 :
(key == 11'b00001000001) ? 46'b0000011100111101100011100000111001111011000111 :
(key == 11'b00001000010) ? 46'b0000011100011110101001100000111000111101010011 :
(key == 11'b00001000011) ? 46'b0000011011111111110011000000110111111111100110 :
(key == 11'b00001000100) ? 46'b0000011011100000111110000000110111000001111100 :
(key == 11'b00001000101) ? 46'b0000011011000010001100000000110110000100011000 :
(key == 11'b00001000110) ? 46'b0000011010100011011101000000110101000110111010 :
(key == 11'b00001000111) ? 46'b0000011010000100110000000000110100001001100000 :
(key == 11'b00001001000) ? 46'b0000011001100110000110100000110011001100001101 :
(key == 11'b00001001001) ? 46'b0000011001000111100000000000110010001111000000 :
(key == 11'b00001001010) ? 46'b0000011000101000111011100000110001010001110111 :
(key == 11'b00001001011) ? 46'b0000011000001010011001100000110000010100110011 :
(key == 11'b00001001100) ? 46'b0000010111101011111010000000101111010111110100 :
(key == 11'b00001001101) ? 46'b0000010111001101011110000000101110011010111100 :
(key == 11'b00001001110) ? 46'b0000010110101111000100000000101101011110001000 :
(key == 11'b00001001111) ? 46'b0000010110010000101101100000101100100001011011 :
(key == 11'b00001010000) ? 46'b0000010101110010011001000000101011100100110010 :
(key == 11'b00001010001) ? 46'b0000010101010100000111000000101010101000001110 :
(key == 11'b00001010010) ? 46'b0000010100110101111000000000101001101011110000 :
(key == 11'b00001010011) ? 46'b0000010100010111101011100000101000101111010111 :
(key == 11'b00001010100) ? 46'b0000010011111001100001000000100111110011000010 :
(key == 11'b00001010101) ? 46'b0000010011011011011010000000100110110110110100 :
(key == 11'b00001010110) ? 46'b0000010010111101010101000000100101111010101010 :
(key == 11'b00001010111) ? 46'b0000010010011111010011000000100100111110100110 :
(key == 11'b00001011000) ? 46'b0000010010000001010100000000100100000010101000 :
(key == 11'b00001011001) ? 46'b0000010001100011010110100000100011000110101101 :
(key == 11'b00001011010) ? 46'b0000010001000101011100000000100010001010111000 :
(key == 11'b00001011011) ? 46'b0000010000100111100100000000100001001111001000 :
(key == 11'b00001011100) ? 46'b0000010000001001101111000000100000010011011110 :
(key == 11'b00001011101) ? 46'b0000001111101011111100000000011111010111111000 :
(key == 11'b00001011110) ? 46'b0000001111001110001100100000011110011100011001 :
(key == 11'b00001011111) ? 46'b0000001110110000011111000000011101100000111110 :
(key == 11'b00001100000) ? 46'b0000001110010010110100000000011100100101101000 :
(key == 11'b00001100001) ? 46'b0000001101110101001011100000011011101010010111 :
(key == 11'b00001100010) ? 46'b0000001101010111100101000000011010101111001010 :
(key == 11'b00001100011) ? 46'b0000001100111010000010000000011001110100000100 :
(key == 11'b00001100100) ? 46'b0000001100011100100001000000011000111001000010 :
(key == 11'b00001100101) ? 46'b0000001011111111000011000000010111111110000110 :
(key == 11'b00001100110) ? 46'b0000001011100001100111000000010111000011001110 :
(key == 11'b00001100111) ? 46'b0000001011000100001101100000010110001000011011 :
(key == 11'b00001101000) ? 46'b0000001010100110110110100000010101001101101101 :
(key == 11'b00001101001) ? 46'b0000001010001001100010100000010100010011000101 :
(key == 11'b00001101010) ? 46'b0000001001101100010000100000010011011000100001 :
(key == 11'b00001101011) ? 46'b0000001001001111000001000000010010011110000010 :
(key == 11'b00001101100) ? 46'b0000001000110001110100000000010001100011101000 :
(key == 11'b00001101101) ? 46'b0000001000010100101010000000010000101001010100 :
(key == 11'b00001101110) ? 46'b0000000111110111100010000000001111101111000100 :
(key == 11'b00001101111) ? 46'b0000000111011010011100000000001110110100111000 :
(key == 11'b00001110000) ? 46'b0000000110111101011001100000001101111010110011 :
(key == 11'b00001110001) ? 46'b0000000110100000011001000000001101000000110010 :
(key == 11'b00001110010) ? 46'b0000000110000011011010100000001100000110110101 :
(key == 11'b00001110011) ? 46'b0000000101100110011111000000001011001100111110 :
(key == 11'b00001110100) ? 46'b0000000101001001100101100000001010010011001011 :
(key == 11'b00001110101) ? 46'b0000000100101100101110100000001001011001011101 :
(key == 11'b00001110110) ? 46'b0000000100001111111010000000001000011111110100 :
(key == 11'b00001110111) ? 46'b0000000011110011001000000000000111100110010000 :
(key == 11'b00001111000) ? 46'b0000000011010110011000100000000110101100110001 :
(key == 11'b00001111001) ? 46'b0000000010111001101011100000000101110011010111 :
(key == 11'b00001111010) ? 46'b0000000010011101000000100000000100111010000001 :
(key == 11'b00001111011) ? 46'b0000000010000000011000000000000100000000110000 :
(key == 11'b00001111100) ? 46'b0000000001100011110010100000000011000111100101 :
(key == 11'b00001111101) ? 46'b0000000001000111001110100000000010001110011101 :
(key == 11'b00001111110) ? 46'b0000000000101010101101100000000001010101011011 :
(key == 11'b00001111111) ? 46'b0000000000001110001111000000000000011100011110 :
(key == 11'b00010000000) ? 46'b1111111111100011100101111111111111000111001011 :
(key == 11'b00010000001) ? 46'b1111111110101010110001011111111101010101100010 :
(key == 11'b00010000010) ? 46'b1111111101110010000000111111111011100100000001 :
(key == 11'b00010000011) ? 46'b1111111100111001010110011111111001110010101100 :
(key == 11'b00010000100) ? 46'b1111111100000000110000111111111000000001100001 :
(key == 11'b00010000101) ? 46'b1111111011001000001111011111110110010000011110 :
(key == 11'b00010000110) ? 46'b1111111010001111110010111111110100011111100101 :
(key == 11'b00010000111) ? 46'b1111111001010111011010011111110010101110110100 :
(key == 11'b00010001000) ? 46'b1111111000011111000111011111110000111110001110 :
(key == 11'b00010001001) ? 46'b1111110111100110111001011111101111001101110010 :
(key == 11'b00010001010) ? 46'b1111110110101110101111011111101101011101011110 :
(key == 11'b00010001011) ? 46'b1111110101110110101001011111101011101101010010 :
(key == 11'b00010001100) ? 46'b1111110100111110101001011111101001111101010010 :
(key == 11'b00010001101) ? 46'b1111110100000110101100011111101000001101011000 :
(key == 11'b00010001110) ? 46'b1111110011001110110100111111100110011101101001 :
(key == 11'b00010001111) ? 46'b1111110010010111000010111111100100101110000101 :
(key == 11'b00010010000) ? 46'b1111110001011111010011111111100010111110100111 :
(key == 11'b00010010001) ? 46'b1111110000100111101010011111100001001111010100 :
(key == 11'b00010010010) ? 46'b1111101111110000000100111111011111100000001001 :
(key == 11'b00010010011) ? 46'b1111101110111000100100011111011101110001001000 :
(key == 11'b00010010100) ? 46'b1111101110000001001000011111011100000010010000 :
(key == 11'b00010010101) ? 46'b1111101101001001110000111111011010010011100001 :
(key == 11'b00010010110) ? 46'b1111101100010010011101011111011000100100111010 :
(key == 11'b00010010111) ? 46'b1111101011011011001110111111010110110110011101 :
(key == 11'b00010011000) ? 46'b1111101010100100000100011111010101001000001000 :
(key == 11'b00010011001) ? 46'b1111101001101100111110111111010011011001111101 :
(key == 11'b00010011010) ? 46'b1111101000110101111110011111010001101011111100 :
(key == 11'b00010011011) ? 46'b1111100111111111000010011111001111111110000100 :
(key == 11'b00010011100) ? 46'b1111100111001000001010011111001110010000010100 :
(key == 11'b00010011101) ? 46'b1111100110010001010111011111001100100010101110 :
(key == 11'b00010011110) ? 46'b1111100101011010100111011111001010110101001110 :
(key == 11'b00010011111) ? 46'b1111100100100011111100011111001001000111111000 :
(key == 11'b00010100000) ? 46'b1111100011101101010110111111000111011010101101 :
(key == 11'b00010100001) ? 46'b1111100010110110110101011111000101101101101010 :
(key == 11'b00010100010) ? 46'b1111100010000000010111011111000100000000101110 :
(key == 11'b00010100011) ? 46'b1111100001001001111101011111000010010011111010 :
(key == 11'b00010100100) ? 46'b1111100000010011101001011111000000100111010010 :
(key == 11'b00010100101) ? 46'b1111011111011101011000111110111110111010110001 :
(key == 11'b00010100110) ? 46'b1111011110100111001100111110111101001110011001 :
(key == 11'b00010100111) ? 46'b1111011101110001000101011110111011100010001010 :
(key == 11'b00010101000) ? 46'b1111011100111011000010011110111001110110000100 :
(key == 11'b00010101001) ? 46'b1111011100000101000011011110111000001010000110 :
(key == 11'b00010101010) ? 46'b1111011011001111001001011110110110011110010010 :
(key == 11'b00010101011) ? 46'b1111011010011001010010111110110100110010100101 :
(key == 11'b00010101100) ? 46'b1111011001100011100001011110110011000111000010 :
(key == 11'b00010101101) ? 46'b1111011000101101110011011110110001011011100110 :
(key == 11'b00010101110) ? 46'b1111010111111000001010011110101111110000010100 :
(key == 11'b00010101111) ? 46'b1111010111000010100100011110101110000101001000 :
(key == 11'b00010110000) ? 46'b1111010110001101000100111110101100011010001001 :
(key == 11'b00010110001) ? 46'b1111010101010111101000011110101010101111010000 :
(key == 11'b00010110010) ? 46'b1111010100100010001111111110101001000100011111 :
(key == 11'b00010110011) ? 46'b1111010011101100111100011110100111011001111000 :
(key == 11'b00010110100) ? 46'b1111010010110111101100111110100101101111011001 :
(key == 11'b00010110101) ? 46'b1111010010000010100001011110100100000101000010 :
(key == 11'b00010110110) ? 46'b1111010001001101011010011110100010011010110100 :
(key == 11'b00010110111) ? 46'b1111010000011000010111111110100000110000101111 :
(key == 11'b00010111000) ? 46'b1111001111100011011001011110011111000110110010 :
(key == 11'b00010111001) ? 46'b1111001110101110011110111110011101011100111101 :
(key == 11'b00010111010) ? 46'b1111001101111001100111011110011011110011001110 :
(key == 11'b00010111011) ? 46'b1111001101000100110101011110011010001001101010 :
(key == 11'b00010111100) ? 46'b1111001100010000001000111110011000100000010001 :
(key == 11'b00010111101) ? 46'b1111001011011011011111011110010110110110111110 :
(key == 11'b00010111110) ? 46'b1111001010100110111001011110010101001101110010 :
(key == 11'b00010111111) ? 46'b1111001001110010010110111110010011100100101101 :
(key == 11'b00011000000) ? 46'b1111001000111101111010011110010001111011110100 :
(key == 11'b00011000001) ? 46'b1111001000001001100000011110010000010011000000 :
(key == 11'b00011000010) ? 46'b1111000111010101001011111110001110101010010111 :
(key == 11'b00011000011) ? 46'b1111000110100000111011011110001101000001110110 :
(key == 11'b00011000100) ? 46'b1111000101101100101110011110001011011001011100 :
(key == 11'b00011000101) ? 46'b1111000100111000100101011110001001110001001010 :
(key == 11'b00011000110) ? 46'b1111000100000100100001011110001000001001000010 :
(key == 11'b00011000111) ? 46'b1111000011010000100000111110000110100001000001 :
(key == 11'b00011001000) ? 46'b1111000010011100100100111110000100111001001001 :
(key == 11'b00011001001) ? 46'b1111000001101000101011111110000011010001010111 :
(key == 11'b00011001010) ? 46'b1111000000110100110111011110000001101001101110 :
(key == 11'b00011001011) ? 46'b1111000000000001000111011110000000000010001110 :
(key == 11'b00011001100) ? 46'b1110111111001101011011111101111110011010110111 :
(key == 11'b00011001101) ? 46'b1110111110011001110011011101111100110011100110 :
(key == 11'b00011001110) ? 46'b1110111101100110001110011101111011001100011100 :
(key == 11'b00011001111) ? 46'b1110111100110010101111011101111001100101011110 :
(key == 11'b00011010000) ? 46'b1110111011111111010011011101110111111110100110 :
(key == 11'b00011010001) ? 46'b1110111011001011111010011101110110010111110100 :
(key == 11'b00011010010) ? 46'b1110111010011000100110011101110100110001001100 :
(key == 11'b00011010011) ? 46'b1110111001100101010110011101110011001010101100 :
(key == 11'b00011010100) ? 46'b1110111000110010001011011101110001100100010110 :
(key == 11'b00011010101) ? 46'b1110110111111111000011011101101111111110000110 :
(key == 11'b00011010110) ? 46'b1110110111001011111101111101101110010111111011 :
(key == 11'b00011010111) ? 46'b1110110110011000111101011101101100110001111010 :
(key == 11'b00011011000) ? 46'b1110110101100110000010011101101011001100000100 :
(key == 11'b00011011001) ? 46'b1110110100110011001001111101101001100110010011 :
(key == 11'b00011011010) ? 46'b1110110100000000010101011101101000000000101010 :
(key == 11'b00011011011) ? 46'b1110110011001101100100011101100110011011001000 :
(key == 11'b00011011100) ? 46'b1110110010011010110111011101100100110101101110 :
(key == 11'b00011011101) ? 46'b1110110001101000001110111101100011010000011101 :
(key == 11'b00011011110) ? 46'b1110110000110101101011011101100001101011010110 :
(key == 11'b00011011111) ? 46'b1110110000000011001010011101100000000110010100 :
(key == 11'b00011100000) ? 46'b1110101111010000101100011101011110100001011000 :
(key == 11'b00011100001) ? 46'b1110101110011110010011011101011100111100100110 :
(key == 11'b00011100010) ? 46'b1110101101101011111110011101011011010111111100 :
(key == 11'b00011100011) ? 46'b1110101100111001101100111101011001110011011001 :
(key == 11'b00011100100) ? 46'b1110101100000111011111011101011000001110111110 :
(key == 11'b00011100101) ? 46'b1110101011010101010110011101010110101010101100 :
(key == 11'b00011100110) ? 46'b1110101010100011010000011101010101000110100000 :
(key == 11'b00011100111) ? 46'b1110101001110001001101111101010011100010011011 :
(key == 11'b00011101000) ? 46'b1110101000111111001111111101010001111110011111 :
(key == 11'b00011101001) ? 46'b1110101000001101010101011101010000011010101010 :
(key == 11'b00011101010) ? 46'b1110100111011011011111011101001110110110111110 :
(key == 11'b00011101011) ? 46'b1110100110101001101011011101001101010011010110 :
(key == 11'b00011101100) ? 46'b1110100101110111111101011101001011101111111010 :
(key == 11'b00011101101) ? 46'b1110100101000110010001011101001010001100100010 :
(key == 11'b00011101110) ? 46'b1110100100010100101010011101001000101001010100 :
(key == 11'b00011101111) ? 46'b1110100011100011000111011101000111000110001110 :
(key == 11'b00011110000) ? 46'b1110100010110001100111011101000101100011001110 :
(key == 11'b00011110001) ? 46'b1110100010000000001011011101000100000000010110 :
(key == 11'b00011110010) ? 46'b1110100001001110110010111101000010011101100101 :
(key == 11'b00011110011) ? 46'b1110100000011101011110011101000000111010111100 :
(key == 11'b00011110100) ? 46'b1110011111101100001101011100111111011000011010 :
(key == 11'b00011110101) ? 46'b1110011110111010111111111100111101110101111111 :
(key == 11'b00011110110) ? 46'b1110011110001001110111011100111100010011101110 :
(key == 11'b00011110111) ? 46'b1110011101011000110000011100111010110001100000 :
(key == 11'b00011111000) ? 46'b1110011100100111101110011100111001001111011100 :
(key == 11'b00011111001) ? 46'b1110011011110110110000011100110111101101100000 :
(key == 11'b00011111010) ? 46'b1110011011000101110101111100110110001011101011 :
(key == 11'b00011111011) ? 46'b1110011010010100111111011100110100101001111110 :
(key == 11'b00011111100) ? 46'b1110011001100100001011011100110011001000010110 :
(key == 11'b00011111101) ? 46'b1110011000110011011011011100110001100110110110 :
(key == 11'b00011111110) ? 46'b1110011000000010101111111100110000000101011111 :
(key == 11'b00011111111) ? 46'b1110010111010010000111011100101110100100001110 :
(key == 11'b00100000000) ? 46'b1110010110100001100010011100101101000011000100 :
(key == 11'b00100000001) ? 46'b1110010101110001000010011100101011100010000100 :
(key == 11'b00100000010) ? 46'b1110010101000000100101011100101010000001001010 :
(key == 11'b00100000011) ? 46'b1110010100010000001010111100101000100000010101 :
(key == 11'b00100000100) ? 46'b1110010011011111110100011100100110111111101000 :
(key == 11'b00100000101) ? 46'b1110010010101111100001011100100101011111000010 :
(key == 11'b00100000110) ? 46'b1110010001111111010011011100100011111110100110 :
(key == 11'b00100000111) ? 46'b1110010001001111001000011100100010011110010000 :
(key == 11'b00100001000) ? 46'b1110010000011111000000011100100000111110000000 :
(key == 11'b00100001001) ? 46'b1110001111101110111100111100011111011101111001 :
(key == 11'b00100001010) ? 46'b1110001110111110111100011100011101111101111000 :
(key == 11'b00100001011) ? 46'b1110001110001110111110011100011100011101111100 :
(key == 11'b00100001100) ? 46'b1110001101011111000101011100011010111110001010 :
(key == 11'b00100001101) ? 46'b1110001100101111001111011100011001011110011110 :
(key == 11'b00100001110) ? 46'b1110001011111111011101011100010111111110111010 :
(key == 11'b00100001111) ? 46'b1110001011001111101110011100010110011111011100 :
(key == 11'b00100010000) ? 46'b1110001010100000000011011100010101000000000110 :
(key == 11'b00100010001) ? 46'b1110001001110000011011011100010011100000110110 :
(key == 11'b00100010010) ? 46'b1110001001000000110111011100010010000001101110 :
(key == 11'b00100010011) ? 46'b1110001000010001010110011100010000100010101100 :
(key == 11'b00100010100) ? 46'b1110000111100001111001011100001111000011110010 :
(key == 11'b00100010101) ? 46'b1110000110110010011111011100001101100100111110 :
(key == 11'b00100010110) ? 46'b1110000110000011001001011100001100000110010010 :
(key == 11'b00100010111) ? 46'b1110000101010011110111011100001010100111101110 :
(key == 11'b00100011000) ? 46'b1110000100100100100111011100001001001001001110 :
(key == 11'b00100011001) ? 46'b1110000011110101011011011100000111101010110110 :
(key == 11'b00100011010) ? 46'b1110000011000110010011111100000110001100100111 :
(key == 11'b00100011011) ? 46'b1110000010010111001111011100000100101110011110 :
(key == 11'b00100011100) ? 46'b1110000001101000001110011100000011010000011100 :
(key == 11'b00100011101) ? 46'b1110000000111001001111011100000001110010011110 :
(key == 11'b00100011110) ? 46'b1110000000001010010101011100000000010100101010 :
(key == 11'b00100011111) ? 46'b1101111111011011011101111011111110110110111011 :
(key == 11'b00100100000) ? 46'b1101111110101100101010011011111101011001010100 :
(key == 11'b00100100001) ? 46'b1101111101111101111001111011111011111011110011 :
(key == 11'b00100100010) ? 46'b1101111101001111001101011011111010011110011010 :
(key == 11'b00100100011) ? 46'b1101111100100000100100011011111001000001001000 :
(key == 11'b00100100100) ? 46'b1101111011110001111110011011110111100011111100 :
(key == 11'b00100100101) ? 46'b1101111011000011011011111011110110000110110111 :
(key == 11'b00100100110) ? 46'b1101111010010100111100011011110100101001111000 :
(key == 11'b00100100111) ? 46'b1101111001100110100000011011110011001101000000 :
(key == 11'b00100101000) ? 46'b1101111000111000001000011011110001110000010000 :
(key == 11'b00100101001) ? 46'b1101111000001001110011011011110000010011100110 :
(key == 11'b00100101010) ? 46'b1101110111011011100010011011101110110111000100 :
(key == 11'b00100101011) ? 46'b1101110110101101010011011011101101011010100110 :
(key == 11'b00100101100) ? 46'b1101110101111111000111011011101011111110001110 :
(key == 11'b00100101101) ? 46'b1101110101010000111111011011101010100001111110 :
(key == 11'b00100101110) ? 46'b1101110100100010111011011011101001000101110110 :
(key == 11'b00100101111) ? 46'b1101110011110100111010111011100111101001110101 :
(key == 11'b00100110000) ? 46'b1101110011000110111101011011100110001101111010 :
(key == 11'b00100110001) ? 46'b1101110010011001000010111011100100110010000101 :
(key == 11'b00100110010) ? 46'b1101110001101011001100011011100011010110011000 :
(key == 11'b00100110011) ? 46'b1101110000111101011001011011100001111010110010 :
(key == 11'b00100110100) ? 46'b1101110000001111100111011011100000011111001110 :
(key == 11'b00100110101) ? 46'b1101101111100001111010011011011111000011110100 :
(key == 11'b00100110110) ? 46'b1101101110110100010001011011011101101000100010 :
(key == 11'b00100110111) ? 46'b1101101110000110101010011011011100001101010100 :
(key == 11'b00100111000) ? 46'b1101101101011001000111011011011010110010001110 :
(key == 11'b00100111001) ? 46'b1101101100101011100111011011011001010111001110 :
(key == 11'b00100111010) ? 46'b1101101011111110001010011011010111111100010100 :
(key == 11'b00100111011) ? 46'b1101101011010000110001011011010110100001100010 :
(key == 11'b00100111100) ? 46'b1101101010100011011011011011010101000110110110 :
(key == 11'b00100111101) ? 46'b1101101001110110000111011011010011101100001110 :
(key == 11'b00100111110) ? 46'b1101101001001000110111111011010010010001101111 :
(key == 11'b00100111111) ? 46'b1101101000011011101011111011010000110111010111 :
(key == 11'b00101000000) ? 46'b1101100111101110100010011011001111011101000100 :
(key == 11'b00101000001) ? 46'b1101100111000001011100011011001110000010111000 :
(key == 11'b00101000010) ? 46'b1101100110010100011001011011001100101000110010 :
(key == 11'b00101000011) ? 46'b1101100101100111011001111011001011001110110011 :
(key == 11'b00101000100) ? 46'b1101100100111010011100111011001001110100111001 :
(key == 11'b00101000101) ? 46'b1101100100001101100011011011001000011011000110 :
(key == 11'b00101000110) ? 46'b1101100011100000101110011011000111000001011100 :
(key == 11'b00101000111) ? 46'b1101100010110011111011011011000101100111110110 :
(key == 11'b00101001000) ? 46'b1101100010000111001011011011000100001110010110 :
(key == 11'b00101001001) ? 46'b1101100001011010011111011011000010110100111110 :
(key == 11'b00101001010) ? 46'b1101100000101101110110011011000001011011101100 :
(key == 11'b00101001011) ? 46'b1101100000000001001111011011000000000010011110 :
(key == 11'b00101001100) ? 46'b1101011111010100101100111010111110101001011001 :
(key == 11'b00101001101) ? 46'b1101011110101000001101011010111101010000011010 :
(key == 11'b00101001110) ? 46'b1101011101111011110000011010111011110111100000 :
(key == 11'b00101001111) ? 46'b1101011101001111010110011010111010011110101100 :
(key == 11'b00101010000) ? 46'b1101011100100011000000011010111001000110000000 :
(key == 11'b00101010001) ? 46'b1101011011110110101100111010110111101101011001 :
(key == 11'b00101010010) ? 46'b1101011011001010011100111010110110010100111001 :
(key == 11'b00101010011) ? 46'b1101011010011110001111011010110100111100011110 :
(key == 11'b00101010100) ? 46'b1101011001110010000101111010110011100100001011 :
(key == 11'b00101010101) ? 46'b1101011001000101111110111010110010001011111101 :
(key == 11'b00101010110) ? 46'b1101011000011001111010111010110000110011110101 :
(key == 11'b00101010111) ? 46'b1101010111101101111011011010101111011011110110 :
(key == 11'b00101011000) ? 46'b1101010111000001111101011010101110000011111010 :
(key == 11'b00101011001) ? 46'b1101010110010110000010011010101100101100000100 :
(key == 11'b00101011010) ? 46'b1101010101101010001011011010101011010100010110 :
(key == 11'b00101011011) ? 46'b1101010100111110010110111010101001111100101101 :
(key == 11'b00101011100) ? 46'b1101010100010010100100111010101000100101001001 :
(key == 11'b00101011101) ? 46'b1101010011100110110111011010100111001101101110 :
(key == 11'b00101011110) ? 46'b1101010010111011001100011010100101110110011000 :
(key == 11'b00101011111) ? 46'b1101010010001111100011111010100100011111000111 :
(key == 11'b00101100000) ? 46'b1101010001100011111111011010100011000111111110 :
(key == 11'b00101100001) ? 46'b1101010000111000011101011010100001110000111010 :
(key == 11'b00101100010) ? 46'b1101010000001100111101111010100000011001111011 :
(key == 11'b00101100011) ? 46'b1101001111100001100010011010011111000011000100 :
(key == 11'b00101100100) ? 46'b1101001110110110001001011010011101101100010010 :
(key == 11'b00101100101) ? 46'b1101001110001010110010111010011100010101100101 :
(key == 11'b00101100110) ? 46'b1101001101011111011111011010011010111110111110 :
(key == 11'b00101100111) ? 46'b1101001100110100010000011010011001101000100000 :
(key == 11'b00101101000) ? 46'b1101001100001001000011011010011000010010000110 :
(key == 11'b00101101001) ? 46'b1101001011011101111001011010010110111011110010 :
(key == 11'b00101101010) ? 46'b1101001010110010110010111010010101100101100101 :
(key == 11'b00101101011) ? 46'b1101001010000111101110011010010100001111011100 :
(key == 11'b00101101100) ? 46'b1101001001011100101101011010010010111001011010 :
(key == 11'b00101101101) ? 46'b1101001000110001101111111010010001100011011111 :
(key == 11'b00101101110) ? 46'b1101001000000110110100011010010000001101101000 :
(key == 11'b00101101111) ? 46'b1101000111011011111100011010001110110111111000 :
(key == 11'b00101110000) ? 46'b1101000110110001000111011010001101100010001110 :
(key == 11'b00101110001) ? 46'b1101000110000110010101011010001100001100101010 :
(key == 11'b00101110010) ? 46'b1101000101011011100110011010001010110111001100 :
(key == 11'b00101110011) ? 46'b1101000100110000111010011010001001100001110100 :
(key == 11'b00101110100) ? 46'b1101000100000110010000011010001000001100100000 :
(key == 11'b00101110101) ? 46'b1101000011011011101001111010000110110111010011 :
(key == 11'b00101110110) ? 46'b1101000010110001000110011010000101100010001100 :
(key == 11'b00101110111) ? 46'b1101000010000110100101011010000100001101001010 :
(key == 11'b00101111000) ? 46'b1101000001011100001000011010000010111000010000 :
(key == 11'b00101111001) ? 46'b1101000000110001101101011010000001100011011010 :
(key == 11'b00101111010) ? 46'b1101000000000111010110011010000000001110101100 :
(key == 11'b00101111011) ? 46'b1100111111011101000000011001111110111010000000 :
(key == 11'b00101111100) ? 46'b1100111110110010101110011001111101100101011100 :
(key == 11'b00101111101) ? 46'b1100111110001000011111011001111100010000111110 :
(key == 11'b00101111110) ? 46'b1100111101011110010011011001111010111100100110 :
(key == 11'b00101111111) ? 46'b1100111100110100001001011001111001101000010010 :
(key == 11'b00110000000) ? 46'b1100111100001010000011011001111000010100000110 :
(key == 11'b00110000001) ? 46'b1100111011011111111111111001110110111111111111 :
(key == 11'b00110000010) ? 46'b1100111010110101111111011001110101101011111110 :
(key == 11'b00110000011) ? 46'b1100111010001100000001011001110100011000000010 :
(key == 11'b00110000100) ? 46'b1100111001100010000101111001110011000100001011 :
(key == 11'b00110000101) ? 46'b1100111000111000001110011001110001110000011100 :
(key == 11'b00110000110) ? 46'b1100111000001110010111111001110000011100101111 :
(key == 11'b00110000111) ? 46'b1100110111100100100101011001101111001001001010 :
(key == 11'b00110001000) ? 46'b1100110110111010110101111001101101110101101011 :
(key == 11'b00110001001) ? 46'b1100110110010001001001011001101100100010010010 :
(key == 11'b00110001010) ? 46'b1100110101100111011111011001101011001110111110 :
(key == 11'b00110001011) ? 46'b1100110100111101110111011001101001111011101110 :
(key == 11'b00110001100) ? 46'b1100110100010100010010111001101000101000100101 :
(key == 11'b00110001101) ? 46'b1100110011101010110001011001100111010101100010 :
(key == 11'b00110001110) ? 46'b1100110011000001010010011001100110000010100100 :
(key == 11'b00110001111) ? 46'b1100110010010111110110011001100100101111101100 :
(key == 11'b00110010000) ? 46'b1100110001101110011101011001100011011100111010 :
(key == 11'b00110010001) ? 46'b1100110001000101000110111001100010001010001101 :
(key == 11'b00110010010) ? 46'b1100110000011011110011011001100000110111100110 :
(key == 11'b00110010011) ? 46'b1100101111110010100011011001011111100101000110 :
(key == 11'b00110010100) ? 46'b1100101111001001010100011001011110010010101000 :
(key == 11'b00110010101) ? 46'b1100101110100000001001011001011101000000010010 :
(key == 11'b00110010110) ? 46'b1100101101110111000000011001011011101110000000 :
(key == 11'b00110010111) ? 46'b1100101101001101111010011001011010011011110100 :
(key == 11'b00110011000) ? 46'b1100101100100100110111011001011001001001101110 :
(key == 11'b00110011001) ? 46'b1100101011111011110110111001010111110111101101 :
(key == 11'b00110011010) ? 46'b1100101011010010111001011001010110100101110010 :
(key == 11'b00110011011) ? 46'b1100101010101001111110011001010101010011111100 :
(key == 11'b00110011100) ? 46'b1100101010000001000110011001010100000010001100 :
(key == 11'b00110011101) ? 46'b1100101001011000010000111001010010110000100001 :
(key == 11'b00110011110) ? 46'b1100101000101111011110111001010001011110111101 :
(key == 11'b00110011111) ? 46'b1100101000000110101110011001010000001101011100 :
(key == 11'b00110100000) ? 46'b1100100111011110000001011001001110111100000010 :
(key == 11'b00110100001) ? 46'b1100100110110101010111011001001101101010101110 :
(key == 11'b00110100010) ? 46'b1100100110001100101110111001001100011001011101 :
(key == 11'b00110100011) ? 46'b1100100101100100001010011001001011001000010100 :
(key == 11'b00110100100) ? 46'b1100100100111011100111011001001001110111001110 :
(key == 11'b00110100101) ? 46'b1100100100010011001000011001001000100110010000 :
(key == 11'b00110100110) ? 46'b1100100011101010101011011001000111010101010110 :
(key == 11'b00110100111) ? 46'b1100100011000010010001011001000110000100100010 :
(key == 11'b00110101000) ? 46'b1100100010011001111001011001000100110011110010 :
(key == 11'b00110101001) ? 46'b1100100001110001100100011001000011100011001000 :
(key == 11'b00110101010) ? 46'b1100100001001001010001011001000010010010100010 :
(key == 11'b00110101011) ? 46'b1100100000100001000001111001000001000010000011 :
(key == 11'b00110101100) ? 46'b1100011111111000110101011000111111110001101010 :
(key == 11'b00110101101) ? 46'b1100011111010000101010011000111110100001010100 :
(key == 11'b00110101110) ? 46'b1100011110101000100011011000111101010001000110 :
(key == 11'b00110101111) ? 46'b1100011110000000011110011000111100000000111100 :
(key == 11'b00110110000) ? 46'b1100011101011000011011011000111010110000110110 :
(key == 11'b00110110001) ? 46'b1100011100110000011100011000111001100000111000 :
(key == 11'b00110110010) ? 46'b1100011100001000011110111000111000010000111101 :
(key == 11'b00110110011) ? 46'b1100011011100000100101011000110111000001001010 :
(key == 11'b00110110100) ? 46'b1100011010111000101100011000110101110001011000 :
(key == 11'b00110110101) ? 46'b1100011010010000110110111000110100100001101101 :
(key == 11'b00110110110) ? 46'b1100011001101001000100011000110011010010001000 :
(key == 11'b00110110111) ? 46'b1100011001000001010100011000110010000010101000 :
(key == 11'b00110111000) ? 46'b1100011000011001100110111000110000110011001101 :
(key == 11'b00110111001) ? 46'b1100010111110001111100011000101111100011111000 :
(key == 11'b00110111010) ? 46'b1100010111001010010100011000101110010100101000 :
(key == 11'b00110111011) ? 46'b1100010110100010101110111000101101000101011101 :
(key == 11'b00110111100) ? 46'b1100010101111011001011011000101011110110010110 :
(key == 11'b00110111101) ? 46'b1100010101010011101011011000101010100111010110 :
(key == 11'b00110111110) ? 46'b1100010100101100001101011000101001011000011010 :
(key == 11'b00110111111) ? 46'b1100010100000100110001011000101000001001100010 :
(key == 11'b00111000000) ? 46'b1100010011011101011000111000100110111010110001 :
(key == 11'b00111000001) ? 46'b1100010010110110000011011000100101101100000110 :
(key == 11'b00111000010) ? 46'b1100010010001110101111011000100100011101011110 :
(key == 11'b00111000011) ? 46'b1100010001100111011110011000100011001110111100 :
(key == 11'b00111000100) ? 46'b1100010001000000010000011000100010000000100000 :
(key == 11'b00111000101) ? 46'b1100010000011001000011011000100000110010000110 :
(key == 11'b00111000110) ? 46'b1100001111110001111010011000011111100011110100 :
(key == 11'b00111000111) ? 46'b1100001111001010110100011000011110010101101000 :
(key == 11'b00111001000) ? 46'b1100001110100011101111011000011101000111011110 :
(key == 11'b00111001001) ? 46'b1100001101111100101101011000011011111001011010 :
(key == 11'b00111001010) ? 46'b1100001101010101101110011000011010101011011100 :
(key == 11'b00111001011) ? 46'b1100001100101110110010011000011001011101100100 :
(key == 11'b00111001100) ? 46'b1100001100000111110111011000011000001111101110 :
(key == 11'b00111001101) ? 46'b1100001011100000111111011000010111000001111110 :
(key == 11'b00111001110) ? 46'b1100001010111010001010011000010101110100010100 :
(key == 11'b00111001111) ? 46'b1100001010010011011000011000010100100110110000 :
(key == 11'b00111010000) ? 46'b1100001001101100101000011000010011011001010000 :
(key == 11'b00111010001) ? 46'b1100001001000101111010011000010010001011110100 :
(key == 11'b00111010010) ? 46'b1100001000011111001111011000010000111110011110 :
(key == 11'b00111010011) ? 46'b1100000111111000100111011000001111110001001110 :
(key == 11'b00111010100) ? 46'b1100000111010001111111111000001110100011111111 :
(key == 11'b00111010101) ? 46'b1100000110101011011100011000001101010110111000 :
(key == 11'b00111010110) ? 46'b1100000110000100111011011000001100001001110110 :
(key == 11'b00111010111) ? 46'b1100000101011110011100111000001010111100111001 :
(key == 11'b00111011000) ? 46'b1100000100111000000000011000001001110000000000 :
(key == 11'b00111011001) ? 46'b1100000100010001100110011000001000100011001100 :
(key == 11'b00111011010) ? 46'b1100000011101011001110111000000111010110011101 :
(key == 11'b00111011011) ? 46'b1100000011000100111010011000000110001001110100 :
(key == 11'b00111011100) ? 46'b1100000010011110100111011000000100111101001110 :
(key == 11'b00111011101) ? 46'b1100000001111000010111011000000011110000101110 :
(key == 11'b00111011110) ? 46'b1100000001010010001001011000000010100100010010 :
(key == 11'b00111011111) ? 46'b1100000000101011111110111000000001010111111101 :
(key == 11'b00111100000) ? 46'b1100000000000101110101011000000000001011101010 :
(key == 11'b00111100001) ? 46'b1011111111011111110000010111111110111111100000 :
(key == 11'b00111100010) ? 46'b1011111110111001101011010111111101110011010110 :
(key == 11'b00111100011) ? 46'b1011111110010011101010010111111100100111010100 :
(key == 11'b00111100100) ? 46'b1011111101101101101010110111111011011011010101 :
(key == 11'b00111100101) ? 46'b1011111101000111101111010111111010001111011110 :
(key == 11'b00111100110) ? 46'b1011111100100001110100110111111001000011101001 :
(key == 11'b00111100111) ? 46'b1011111011111011111100110111110111110111111001 :
(key == 11'b00111101000) ? 46'b1011111011010110000111110111110110101100001111 :
(key == 11'b00111101001) ? 46'b1011111010110000010101010111110101100000101010 :
(key == 11'b00111101010) ? 46'b1011111010001010100011110111110100010101000111 :
(key == 11'b00111101011) ? 46'b1011111001100100110101010111110011001001101010 :
(key == 11'b00111101100) ? 46'b1011111000111111001001010111110001111110010010 :
(key == 11'b00111101101) ? 46'b1011111000011001100000010111110000110011000000 :
(key == 11'b00111101110) ? 46'b1011110111110011111001010111101111100111110010 :
(key == 11'b00111101111) ? 46'b1011110111001110010100010111101110011100101000 :
(key == 11'b00111110000) ? 46'b1011110110101000110010010111101101010001100100 :
(key == 11'b00111110001) ? 46'b1011110110000011010011010111101100000110100110 :
(key == 11'b00111110010) ? 46'b1011110101011101110101010111101010111011101010 :
(key == 11'b00111110011) ? 46'b1011110100111000011010010111101001110000110100 :
(key == 11'b00111110100) ? 46'b1011110100010011000010010111101000100110000100 :
(key == 11'b00111110101) ? 46'b1011110011101101101011010111100111011011010110 :
(key == 11'b00111110110) ? 46'b1011110011001000010111010111100110010000101110 :
(key == 11'b00111110111) ? 46'b1011110010100011000100010111100101000110001000 :
(key == 11'b00111111000) ? 46'b1011110001111101110101010111100011111011101010 :
(key == 11'b00111111001) ? 46'b1011110001011000101000010111100010110001010000 :
(key == 11'b00111111010) ? 46'b1011110000110011011110010111100001100110111100 :
(key == 11'b00111111011) ? 46'b1011110000001110010101010111100000011100101010 :
(key == 11'b00111111100) ? 46'b1011101111101001001111010111011111010010011110 :
(key == 11'b00111111101) ? 46'b1011101111000100001011010111011110001000010110 :
(key == 11'b00111111110) ? 46'b1011101110011111001001010111011100111110010010 :
(key == 11'b00111111111) ? 46'b1011101101111010001010010111011011110100010100 :
(key == 11'b01000000000) ? 46'b1011101101010101001101110111011010101010011011 :
(key == 11'b01000000001) ? 46'b1011101100110000010011010111011001100000100110 :
(key == 11'b01000000010) ? 46'b1011101100001011011011110111011000010110110111 :
(key == 11'b01000000011) ? 46'b1011101011100110100101110111010111001101001011 :
(key == 11'b01000000100) ? 46'b1011101011000001110010010111010110000011100100 :
(key == 11'b01000000101) ? 46'b1011101010011101000000010111010100111010000000 :
(key == 11'b01000000110) ? 46'b1011101001111000010001010111010011110000100010 :
(key == 11'b01000000111) ? 46'b1011101001010011100100010111010010100111001000 :
(key == 11'b01000001000) ? 46'b1011101000101110111010010111010001011101110100 :
(key == 11'b01000001001) ? 46'b1011101000001010010010010111010000010100100100 :
(key == 11'b01000001010) ? 46'b1011100111100101101100010111001111001011011000 :
(key == 11'b01000001011) ? 46'b1011100111000001001000010111001110000010010000 :
(key == 11'b01000001100) ? 46'b1011100110011100100110010111001100111001001100 :
(key == 11'b01000001101) ? 46'b1011100101111000000111110111001011110000001111 :
(key == 11'b01000001110) ? 46'b1011100101010011101010010111001010100111010100 :
(key == 11'b01000001111) ? 46'b1011100100101111010000010111001001011110100000 :
(key == 11'b01000010000) ? 46'b1011100100001010111000010111001000010101110000 :
(key == 11'b01000010001) ? 46'b1011100011100110100010010111000111001101000100 :
(key == 11'b01000010010) ? 46'b1011100011000010001110010111000110000100011100 :
(key == 11'b01000010011) ? 46'b1011100010011101111101010111000100111011111010 :
(key == 11'b01000010100) ? 46'b1011100001111001101101010111000011110011011010 :
(key == 11'b01000010101) ? 46'b1011100001010101011111110111000010101010111111 :
(key == 11'b01000010110) ? 46'b1011100000110001010101010111000001100010101010 :
(key == 11'b01000010111) ? 46'b1011100000001101001101010111000000011010011010 :
(key == 11'b01000011000) ? 46'b1011011111101001000110010110111111010010001100 :
(key == 11'b01000011001) ? 46'b1011011111000101000001110110111110001010000011 :
(key == 11'b01000011010) ? 46'b1011011110100000111111010110111101000001111110 :
(key == 11'b01000011011) ? 46'b1011011101111101000000010110111011111010000000 :
(key == 11'b01000011100) ? 46'b1011011101011001000010010110111010110010000100 :
(key == 11'b01000011101) ? 46'b1011011100110101000110010110111001101010001100 :
(key == 11'b01000011110) ? 46'b1011011100010001001101110110111000100010011011 :
(key == 11'b01000011111) ? 46'b1011011011101101010110110110110111011010101101 :
(key == 11'b01000100000) ? 46'b1011011011001001100010010110110110010011000100 :
(key == 11'b01000100001) ? 46'b1011011010100101101111010110110101001011011110 :
(key == 11'b01000100010) ? 46'b1011011010000001111110010110110100000011111100 :
(key == 11'b01000100011) ? 46'b1011011001011110010000010110110010111100100000 :
(key == 11'b01000100100) ? 46'b1011011000111010100100110110110001110101001001 :
(key == 11'b01000100101) ? 46'b1011011000010110111010010110110000101101110100 :
(key == 11'b01000100110) ? 46'b1011010111110011010011010110101111100110100110 :
(key == 11'b01000100111) ? 46'b1011010111001111101101010110101110011111011010 :
(key == 11'b01000101000) ? 46'b1011010110101100001010010110101101011000010100 :
(key == 11'b01000101001) ? 46'b1011010110001000101000110110101100010001010001 :
(key == 11'b01000101010) ? 46'b1011010101100101001001110110101011001010010011 :
(key == 11'b01000101011) ? 46'b1011010101000001101101010110101010000011011010 :
(key == 11'b01000101100) ? 46'b1011010100011110010001110110101000111100100011 :
(key == 11'b01000101101) ? 46'b1011010011111010111001010110100111110101110010 :
(key == 11'b01000101110) ? 46'b1011010011010111100010110110100110101111000101 :
(key == 11'b01000101111) ? 46'b1011010010110100001111010110100101101000011110 :
(key == 11'b01000110000) ? 46'b1011010010010000111100110110100100100001111001 :
(key == 11'b01000110001) ? 46'b1011010001101101101100110110100011011011011001 :
(key == 11'b01000110010) ? 46'b1011010001001010011110010110100010010100111100 :
(key == 11'b01000110011) ? 46'b1011010000100111010011010110100001001110100110 :
(key == 11'b01000110100) ? 46'b1011010000000100001001010110100000001000010010 :
(key == 11'b01000110101) ? 46'b1011001111100001000001110110011111000010000011 :
(key == 11'b01000110110) ? 46'b1011001110111101111101010110011101111011111010 :
(key == 11'b01000110111) ? 46'b1011001110011010111001110110011100110101110011 :
(key == 11'b01000111000) ? 46'b1011001101110111111000010110011011101111110000 :
(key == 11'b01000111001) ? 46'b1011001101010100111001010110011010101001110010 :
(key == 11'b01000111010) ? 46'b1011001100110001111100010110011001100011111000 :
(key == 11'b01000111011) ? 46'b1011001100001111000001110110011000011110000011 :
(key == 11'b01000111100) ? 46'b1011001011101100001000010110010111011000010000 :
(key == 11'b01000111101) ? 46'b1011001011001001010010010110010110010010100100 :
(key == 11'b01000111110) ? 46'b1011001010100110011101010110010101001100111010 :
(key == 11'b01000111111) ? 46'b1011001010000011101010110110010100000111010101 :
(key == 11'b01001000000) ? 46'b1011001001100000111011010110010011000001110110 :
(key == 11'b01001000001) ? 46'b1011001000111110001100010110010001111100011000 :
(key == 11'b01001000010) ? 46'b1011001000011011011111010110010000110110111110 :
(key == 11'b01001000011) ? 46'b1011000111111000110101010110001111110001101010 :
(key == 11'b01001000100) ? 46'b1011000111010110001110010110001110101100011100 :
(key == 11'b01001000101) ? 46'b1011000110110011101000010110001101100111010000 :
(key == 11'b01001000110) ? 46'b1011000110010001000100010110001100100010001000 :
(key == 11'b01001000111) ? 46'b1011000101101110100010010110001011011101000100 :
(key == 11'b01001001000) ? 46'b1011000101001100000010010110001010011000000100 :
(key == 11'b01001001001) ? 46'b1011000100101001100100010110001001010011001000 :
(key == 11'b01001001010) ? 46'b1011000100000111001000110110001000001110010001 :
(key == 11'b01001001011) ? 46'b1011000011100100101111010110000111001001011110 :
(key == 11'b01001001100) ? 46'b1011000011000010010111110110000110000100101111 :
(key == 11'b01001001101) ? 46'b1011000010100000000010010110000101000000000100 :
(key == 11'b01001001110) ? 46'b1011000001111101101111010110000011111011011110 :
(key == 11'b01001001111) ? 46'b1011000001011011011110010110000010110110111100 :
(key == 11'b01001010000) ? 46'b1011000000111001001101110110000001110010011011 :
(key == 11'b01001010001) ? 46'b1011000000010111000000010110000000101110000000 :
(key == 11'b01001010010) ? 46'b1010111111110100110101010101111111101001101010 :
(key == 11'b01001010011) ? 46'b1010111111010010101100010101111110100101011000 :
(key == 11'b01001010100) ? 46'b1010111110110000100100110101111101100001001001 :
(key == 11'b01001010101) ? 46'b1010111110001110011111110101111100011100111111 :
(key == 11'b01001010110) ? 46'b1010111101101100011100010101111011011000111000 :
(key == 11'b01001010111) ? 46'b1010111101001010011011010101111010010100110110 :
(key == 11'b01001011000) ? 46'b1010111100101000011100010101111001010000111000 :
(key == 11'b01001011001) ? 46'b1010111100000110011110010101111000001100111100 :
(key == 11'b01001011010) ? 46'b1010111011100100100011010101110111001001000110 :
(key == 11'b01001011011) ? 46'b1010111011000010101010010101110110000101010100 :
(key == 11'b01001011100) ? 46'b1010111010100000110010110101110101000001100101 :
(key == 11'b01001011101) ? 46'b1010111001111110111101010101110011111101111010 :
(key == 11'b01001011110) ? 46'b1010111001011101001010010101110010111010010100 :
(key == 11'b01001011111) ? 46'b1010111000111011011001010101110001110110110010 :
(key == 11'b01001100000) ? 46'b1010111000011001101001010101110000110011010010 :
(key == 11'b01001100001) ? 46'b1010110111110111111100010101101111101111111000 :
(key == 11'b01001100010) ? 46'b1010110111010110010000010101101110101100100000 :
(key == 11'b01001100011) ? 46'b1010110110110100100111010101101101101001001110 :
(key == 11'b01001100100) ? 46'b1010110110010011000000010101101100100110000000 :
(key == 11'b01001100101) ? 46'b1010110101110001011010110101101011100010110101 :
(key == 11'b01001100110) ? 46'b1010110101001111110111010101101010011111101110 :
(key == 11'b01001100111) ? 46'b1010110100101110010101110101101001011100101011 :
(key == 11'b01001101000) ? 46'b1010110100001100110110010101101000011001101100 :
(key == 11'b01001101001) ? 46'b1010110011101011011001010101100111010110110010 :
(key == 11'b01001101010) ? 46'b1010110011001001111101010101100110010011111010 :
(key == 11'b01001101011) ? 46'b1010110010101000100100010101100101010001001000 :
(key == 11'b01001101100) ? 46'b1010110010000111001100010101100100001110011000 :
(key == 11'b01001101101) ? 46'b1010110001100101110110010101100011001011101100 :
(key == 11'b01001101110) ? 46'b1010110001000100100010010101100010001001000100 :
(key == 11'b01001101111) ? 46'b1010110000100011010001010101100001000110100010 :
(key == 11'b01001110000) ? 46'b1010110000000010000001010101100000000100000010 :
(key == 11'b01001110001) ? 46'b1010101111100000110011010101011111000001100110 :
(key == 11'b01001110010) ? 46'b1010101110111111100110010101011101111111001100 :
(key == 11'b01001110011) ? 46'b1010101110011110011101010101011100111100111010 :
(key == 11'b01001110100) ? 46'b1010101101111101010101010101011011111010101010 :
(key == 11'b01001110101) ? 46'b1010101101011100001110010101011010111000011100 :
(key == 11'b01001110110) ? 46'b1010101100111011001010010101011001110110010100 :
(key == 11'b01001110111) ? 46'b1010101100011010000111110101011000110100001111 :
(key == 11'b01001111000) ? 46'b1010101011111001000111010101010111110010001110 :
(key == 11'b01001111001) ? 46'b1010101011011000001000010101010110110000010000 :
(key == 11'b01001111010) ? 46'b1010101010110111001011010101010101101110010110 :
(key == 11'b01001111011) ? 46'b1010101010010110010001010101010100101100100010 :
(key == 11'b01001111100) ? 46'b1010101001110101011000010101010011101010110000 :
(key == 11'b01001111101) ? 46'b1010101001010100100001010101010010101001000010 :
(key == 11'b01001111110) ? 46'b1010101000110011101100010101010001100111011000 :
(key == 11'b01001111111) ? 46'b1010101000010010111001010101010000100101110010 :
(key == 11'b01010000000) ? 46'b1010100111110010000111010101001111100100001110 :
(key == 11'b01010000001) ? 46'b1010100111010001011000110101001110100010110001 :
(key == 11'b01010000010) ? 46'b1010100110110000101010110101001101100001010101 :
(key == 11'b01010000011) ? 46'b1010100110001111111111010101001100011111111110 :
(key == 11'b01010000100) ? 46'b1010100101101111010101010101001011011110101010 :
(key == 11'b01010000101) ? 46'b1010100101001110101101010101001010011101011010 :
(key == 11'b01010000110) ? 46'b1010100100101110000111110101001001011100001111 :
(key == 11'b01010000111) ? 46'b1010100100001101100100010101001000011011001000 :
(key == 11'b01010001000) ? 46'b1010100011101101000010010101000111011010000100 :
(key == 11'b01010001001) ? 46'b1010100011001100100001010101000110011001000010 :
(key == 11'b01010001010) ? 46'b1010100010101100000010010101000101011000000100 :
(key == 11'b01010001011) ? 46'b1010100010001011100110010101000100010111001100 :
(key == 11'b01010001100) ? 46'b1010100001101011001010110101000011010110010101 :
(key == 11'b01010001101) ? 46'b1010100001001010110001110101000010010101100011 :
(key == 11'b01010001110) ? 46'b1010100000101010011011110101000001010100110111 :
(key == 11'b01010001111) ? 46'b1010100000001010000110010101000000010100001100 :
(key == 11'b01010010000) ? 46'b1010011111101001110010010100111111010011100100 :
(key == 11'b01010010001) ? 46'b1010011111001001100000010100111110010011000000 :
(key == 11'b01010010010) ? 46'b1010011110101001010001010100111101010010100010 :
(key == 11'b01010010011) ? 46'b1010011110001001000011010100111100010010000110 :
(key == 11'b01010010100) ? 46'b1010011101101000110111010100111011010001101110 :
(key == 11'b01010010101) ? 46'b1010011101001000101101010100111010010001011010 :
(key == 11'b01010010110) ? 46'b1010011100101000100100110100111001010001001001 :
(key == 11'b01010010111) ? 46'b1010011100001000011110010100111000010000111100 :
(key == 11'b01010011000) ? 46'b1010011011101000011001010100110111010000110010 :
(key == 11'b01010011001) ? 46'b1010011011001000010110010100110110010000101100 :
(key == 11'b01010011010) ? 46'b1010011010101000010110010100110101010000101100 :
(key == 11'b01010011011) ? 46'b1010011010001000010110010100110100010000101100 :
(key == 11'b01010011100) ? 46'b1010011001101000011001010100110011010000110010 :
(key == 11'b01010011101) ? 46'b1010011001001000011101110100110010010000111011 :
(key == 11'b01010011110) ? 46'b1010011000101000100011010100110001010001000110 :
(key == 11'b01010011111) ? 46'b1010011000001000101011010100110000010001010110 :
(key == 11'b01010100000) ? 46'b1010010111101000110101010100101111010001101010 :
(key == 11'b01010100001) ? 46'b1010010111001001000000110100101110010010000001 :
(key == 11'b01010100010) ? 46'b1010010110101001001110010100101101010010011100 :
(key == 11'b01010100011) ? 46'b1010010110001001011101010100101100010010111010 :
(key == 11'b01010100100) ? 46'b1010010101101001101110010100101011010011011100 :
(key == 11'b01010100101) ? 46'b1010010101001010000001010100101010010100000010 :
(key == 11'b01010100110) ? 46'b1010010100101010010101110100101001010100101011 :
(key == 11'b01010100111) ? 46'b1010010100001010101100110100101000010101011001 :
(key == 11'b01010101000) ? 46'b1010010011101011000100010100100111010110001000 :
(key == 11'b01010101001) ? 46'b1010010011001011011101110100100110010110111011 :
(key == 11'b01010101010) ? 46'b1010010010101011111010010100100101010111110100 :
(key == 11'b01010101011) ? 46'b1010010010001100010111010100100100011000101110 :
(key == 11'b01010101100) ? 46'b1010010001101100110111010100100011011001101110 :
(key == 11'b01010101101) ? 46'b1010010001001101010111110100100010011010101111 :
(key == 11'b01010101110) ? 46'b1010010000101101111010010100100001011011110100 :
(key == 11'b01010101111) ? 46'b1010010000001110011111010100100000011100111110 :
(key == 11'b01010110000) ? 46'b1010001111101111000101010100011111011110001010 :
(key == 11'b01010110001) ? 46'b1010001111001111101100110100011110011111011001 :
(key == 11'b01010110010) ? 46'b1010001110110000010110010100011101100000101100 :
(key == 11'b01010110011) ? 46'b1010001110010001000010010100011100100010000100 :
(key == 11'b01010110100) ? 46'b1010001101110001101111010100011011100011011110 :
(key == 11'b01010110101) ? 46'b1010001101010010011111010100011010100100111110 :
(key == 11'b01010110110) ? 46'b1010001100110011001111010100011001100110011110 :
(key == 11'b01010110111) ? 46'b1010001100010100000010010100011000101000000100 :
(key == 11'b01010111000) ? 46'b1010001011110100110111010100010111101001101110 :
(key == 11'b01010111001) ? 46'b1010001011010101101101010100010110101011011010 :
(key == 11'b01010111010) ? 46'b1010001010110110100100010100010101101101001000 :
(key == 11'b01010111011) ? 46'b1010001010010111011101110100010100101110111011 :
(key == 11'b01010111100) ? 46'b1010001001111000011001010100010011110000110010 :
(key == 11'b01010111101) ? 46'b1010001001011001010110010100010010110010101100 :
(key == 11'b01010111110) ? 46'b1010001000111010010100110100010001110100101001 :
(key == 11'b01010111111) ? 46'b1010001000011011010101010100010000110110101010 :
(key == 11'b01011000000) ? 46'b1010000111111100011000010100001111111000110000 :
(key == 11'b01011000001) ? 46'b1010000111011101011011010100001110111010110110 :
(key == 11'b01011000010) ? 46'b1010000110111110100000010100001101111101000000 :
(key == 11'b01011000011) ? 46'b1010000110011111101000010100001100111111010000 :
(key == 11'b01011000100) ? 46'b1010000110000000110001010100001100000001100010 :
(key == 11'b01011000101) ? 46'b1010000101100001111100010100001011000011111000 :
(key == 11'b01011000110) ? 46'b1010000101000011001000010100001010000110010000 :
(key == 11'b01011000111) ? 46'b1010000100100100010110010100001001001000101100 :
(key == 11'b01011001000) ? 46'b1010000100000101100110010100001000001011001100 :
(key == 11'b01011001001) ? 46'b1010000011100110110111010100000111001101101110 :
(key == 11'b01011001010) ? 46'b1010000011001000001010010100000110010000010100 :
(key == 11'b01011001011) ? 46'b1010000010101001011111110100000101010010111111 :
(key == 11'b01011001100) ? 46'b1010000010001010110110010100000100010101101100 :
(key == 11'b01011001101) ? 46'b1010000001101100001110110100000011011000011101 :
(key == 11'b01011001110) ? 46'b1010000001001101101000010100000010011011010000 :
(key == 11'b01011001111) ? 46'b1010000000101111000100010100000001011110001000 :
(key == 11'b01011010000) ? 46'b1010000000010000100010010100000000100001000100 :
(key == 11'b01011010001) ? 46'b1001111111110010000001010011111111100100000010 :
(key == 11'b01011010010) ? 46'b1001111111010011100001010011111110100111000010 :
(key == 11'b01011010011) ? 46'b1001111110110101000011010011111101101010000110 :
(key == 11'b01011010100) ? 46'b1001111110010110100111110011111100101101001111 :
(key == 11'b01011010101) ? 46'b1001111101111000001110010011111011110000011100 :
(key == 11'b01011010110) ? 46'b1001111101011001110101010011111010110011101010 :
(key == 11'b01011010111) ? 46'b1001111100111011011110010011111001110110111100 :
(key == 11'b01011011000) ? 46'b1001111100011101001000010011111000111010010000 :
(key == 11'b01011011001) ? 46'b1001111011111110110101110011110111111101101011 :
(key == 11'b01011011010) ? 46'b1001111011100000100011110011110111000001000111 :
(key == 11'b01011011011) ? 46'b1001111011000010010011010011110110000100100110 :
(key == 11'b01011011100) ? 46'b1001111010100100000101010011110101001000001010 :
(key == 11'b01011011101) ? 46'b1001111010000101111000010011110100001011110000 :
(key == 11'b01011011110) ? 46'b1001111001100111101101010011110011001111011010 :
(key == 11'b01011011111) ? 46'b1001111001001001100010010011110010010011000100 :
(key == 11'b01011100000) ? 46'b1001111000101011011010010011110001010110110100 :
(key == 11'b01011100001) ? 46'b1001111000001101010011010011110000011010100110 :
(key == 11'b01011100010) ? 46'b1001110111101111001111010011101111011110011110 :
(key == 11'b01011100011) ? 46'b1001110111010001001100010011101110100010011000 :
(key == 11'b01011100100) ? 46'b1001110110110011001011010011101101100110010110 :
(key == 11'b01011100101) ? 46'b1001110110010101001011010011101100101010010110 :
(key == 11'b01011100110) ? 46'b1001110101110111001100110011101011101110011001 :
(key == 11'b01011100111) ? 46'b1001110101011001010000010011101010110010100000 :
(key == 11'b01011101000) ? 46'b1001110100111011010101010011101001110110101010 :
(key == 11'b01011101001) ? 46'b1001110100011101011011110011101000111010110111 :
(key == 11'b01011101010) ? 46'b1001110011111111100100010011100111111111001000 :
(key == 11'b01011101011) ? 46'b1001110011100001101101110011100111000011011011 :
(key == 11'b01011101100) ? 46'b1001110011000011111001010011100110000111110010 :
(key == 11'b01011101101) ? 46'b1001110010100110000110010011100101001100001100 :
(key == 11'b01011101110) ? 46'b1001110010001000010100110011100100010000101001 :
(key == 11'b01011101111) ? 46'b1001110001101010100110010011100011010101001100 :
(key == 11'b01011110000) ? 46'b1001110001001100110111010011100010011001101110 :
(key == 11'b01011110001) ? 46'b1001110000101111001011010011100001011110010110 :
(key == 11'b01011110010) ? 46'b1001110000010001100000010011100000100011000000 :
(key == 11'b01011110011) ? 46'b1001101111110011110111110011011111100111101111 :
(key == 11'b01011110100) ? 46'b1001101111010110001111110011011110101100011111 :
(key == 11'b01011110101) ? 46'b1001101110111000101001010011011101110001010010 :
(key == 11'b01011110110) ? 46'b1001101110011011000101010011011100110110001010 :
(key == 11'b01011110111) ? 46'b1001101101111101100010010011011011111011000100 :
(key == 11'b01011111000) ? 46'b1001101101100000000001010011011011000000000010 :
(key == 11'b01011111001) ? 46'b1001101101000010100001010011011010000101000010 :
(key == 11'b01011111010) ? 46'b1001101100100101000011010011011001001010000110 :
(key == 11'b01011111011) ? 46'b1001101100000111100111010011011000001111001110 :
(key == 11'b01011111100) ? 46'b1001101011101010001011110011010111010100010111 :
(key == 11'b01011111101) ? 46'b1001101011001100110010010011010110011001100100 :
(key == 11'b01011111110) ? 46'b1001101010101111011001110011010101011110110011 :
(key == 11'b01011111111) ? 46'b1001101010010010000100010011010100100100001000 :
(key == 11'b01100000000) ? 46'b1001101001110100110000010011010011101001100000 :
(key == 11'b01100000001) ? 46'b1001101001010111011101010011010010101110111010 :
(key == 11'b01100000010) ? 46'b1001101000111010001010110011010001110100010101 :
(key == 11'b01100000011) ? 46'b1001101000011100111010110011010000111001110101 :
(key == 11'b01100000100) ? 46'b1001100111111111101101010011001111111111011010 :
(key == 11'b01100000101) ? 46'b1001100111100010100000010011001111000101000000 :
(key == 11'b01100000110) ? 46'b1001100111000101010100010011001110001010101000 :
(key == 11'b01100000111) ? 46'b1001100110101000001011010011001101010000010110 :
(key == 11'b01100001000) ? 46'b1001100110001011000010110011001100010110000101 :
(key == 11'b01100001001) ? 46'b1001100101101101111100010011001011011011111000 :
(key == 11'b01100001010) ? 46'b1001100101010000110111110011001010100001101111 :
(key == 11'b01100001011) ? 46'b1001100100110011110011110011001001100111100111 :
(key == 11'b01100001100) ? 46'b1001100100010110110010010011001000101101100100 :
(key == 11'b01100001101) ? 46'b1001100011111001110001010011000111110011100010 :
(key == 11'b01100001110) ? 46'b1001100011011100110011010011000110111001100110 :
(key == 11'b01100001111) ? 46'b1001100010111111110101010011000101111111101010 :
(key == 11'b01100010000) ? 46'b1001100010100010111001010011000101000101110010 :
(key == 11'b01100010001) ? 46'b1001100010000101111111110011000100001011111111 :
(key == 11'b01100010010) ? 46'b1001100001101001000111010011000011010010001110 :
(key == 11'b01100010011) ? 46'b1001100001001100001111010011000010011000011110 :
(key == 11'b01100010100) ? 46'b1001100000101111011001010011000001011110110010 :
(key == 11'b01100010101) ? 46'b1001100000010010100101110011000000100101001011 :
(key == 11'b01100010110) ? 46'b1001011111110101110011010010111111101011100110 :
(key == 11'b01100010111) ? 46'b1001011111011001000001110010111110110010000011 :
(key == 11'b01100011000) ? 46'b1001011110111100010010010010111101111000100100 :
(key == 11'b01100011001) ? 46'b1001011110011111100011110010111100111111000111 :
(key == 11'b01100011010) ? 46'b1001011110000010110111110010111100000101101111 :
(key == 11'b01100011011) ? 46'b1001011101100110001101010010111011001100011010 :
(key == 11'b01100011100) ? 46'b1001011101001001100011010010111010010011000110 :
(key == 11'b01100011101) ? 46'b1001011100101100111011010010111001011001110110 :
(key == 11'b01100011110) ? 46'b1001011100010000010100010010111000100000101000 :
(key == 11'b01100011111) ? 46'b1001011011110011110000010010110111100111100000 :
(key == 11'b01100100000) ? 46'b1001011011010111001101010010110110101110011010 :
(key == 11'b01100100001) ? 46'b1001011010111010101010010010110101110101010100 :
(key == 11'b01100100010) ? 46'b1001011010011110001010010010110100111100010100 :
(key == 11'b01100100011) ? 46'b1001011010000001101011010010110100000011010110 :
(key == 11'b01100100100) ? 46'b1001011001100101001101110010110011001010011011 :
(key == 11'b01100100101) ? 46'b1001011001001000110001010010110010010001100010 :
(key == 11'b01100100110) ? 46'b1001011000101100010111010010110001011000101110 :
(key == 11'b01100100111) ? 46'b1001011000001111111110010010110000011111111100 :
(key == 11'b01100101000) ? 46'b1001010111110011100110010010101111100111001100 :
(key == 11'b01100101001) ? 46'b1001010111010111010001010010101110101110100010 :
(key == 11'b01100101010) ? 46'b1001010110111010111100010010101101110101111000 :
(key == 11'b01100101011) ? 46'b1001010110011110101001010010101100111101010010 :
(key == 11'b01100101100) ? 46'b1001010110000010011000010010101100000100110000 :
(key == 11'b01100101101) ? 46'b1001010101100110000111110010101011001100001111 :
(key == 11'b01100101110) ? 46'b1001010101001001111000010010101010010011110000 :
(key == 11'b01100101111) ? 46'b1001010100101101101011110010101001011011010111 :
(key == 11'b01100110000) ? 46'b1001010100010001100000010010101000100011000000 :
(key == 11'b01100110001) ? 46'b1001010011110101010101110010100111101010101011 :
(key == 11'b01100110010) ? 46'b1001010011011001001101010010100110110010011010 :
(key == 11'b01100110011) ? 46'b1001010010111101000101110010100101111010001011 :
(key == 11'b01100110100) ? 46'b1001010010100001000000010010100101000010000000 :
(key == 11'b01100110101) ? 46'b1001010010000100111011110010100100001001110111 :
(key == 11'b01100110110) ? 46'b1001010001101000111001010010100011010001110010 :
(key == 11'b01100110111) ? 46'b1001010001001100110111010010100010011001101110 :
(key == 11'b01100111000) ? 46'b1001010000110000110111010010100001100001101110 :
(key == 11'b01100111001) ? 46'b1001010000010100111000010010100000101001110000 :
(key == 11'b01100111010) ? 46'b1001001111111000111011010010011111110001110110 :
(key == 11'b01100111011) ? 46'b1001001111011100111111010010011110111001111110 :
(key == 11'b01100111100) ? 46'b1001001111000001000101110010011110000010001011 :
(key == 11'b01100111101) ? 46'b1001001110100101001101010010011101001010011010 :
(key == 11'b01100111110) ? 46'b1001001110001001010110010010011100010010101100 :
(key == 11'b01100111111) ? 46'b1001001101101101100000010010011011011011000000 :
(key == 11'b01101000000) ? 46'b1001001101010001101100010010011010100011011000 :
(key == 11'b01101000001) ? 46'b1001001100110101111001010010011001101011110010 :
(key == 11'b01101000010) ? 46'b1001001100011010000111110010011000110100001111 :
(key == 11'b01101000011) ? 46'b1001001011111110010111010010010111111100101110 :
(key == 11'b01101000100) ? 46'b1001001011100010101000010010010111000101010000 :
(key == 11'b01101000101) ? 46'b1001001011000110111010110010010110001101110101 :
(key == 11'b01101000110) ? 46'b1001001010101011001111010010010101010110011110 :
(key == 11'b01101000111) ? 46'b1001001010001111100101010010010100011111001010 :
(key == 11'b01101001000) ? 46'b1001001001110011111100010010010011100111111000 :
(key == 11'b01101001001) ? 46'b1001001001011000010100010010010010110000101000 :
(key == 11'b01101001010) ? 46'b1001001000111100101110010010010001111001011100 :
(key == 11'b01101001011) ? 46'b1001001000100001001001010010010001000010010010 :
(key == 11'b01101001100) ? 46'b1001001000000101100110110010010000001011001101 :
(key == 11'b01101001101) ? 46'b1001000111101010000101010010001111010100001010 :
(key == 11'b01101001110) ? 46'b1001000111001110100100010010001110011101001000 :
(key == 11'b01101001111) ? 46'b1001000110110011000101010010001101100110001010 :
(key == 11'b01101010000) ? 46'b1001000110010111100110010010001100101111001100 :
(key == 11'b01101010001) ? 46'b1001000101111100001010110010001011111000010101 :
(key == 11'b01101010010) ? 46'b1001000101100000101111110010001011000001011111 :
(key == 11'b01101010011) ? 46'b1001000101000101010111010010001010001010101110 :
(key == 11'b01101010100) ? 46'b1001000100101001111110010010001001010011111100 :
(key == 11'b01101010101) ? 46'b1001000100001110101000010010001000011101010000 :
(key == 11'b01101010110) ? 46'b1001000011110011010010110010000111100110100101 :
(key == 11'b01101010111) ? 46'b1001000011010111111111010010000110101111111110 :
(key == 11'b01101011000) ? 46'b1001000010111100101100010010000101111001011000 :
(key == 11'b01101011001) ? 46'b1001000010100001011100010010000101000010111000 :
(key == 11'b01101011010) ? 46'b1001000010000110001100010010000100001100011000 :
(key == 11'b01101011011) ? 46'b1001000001101010111110010010000011010101111100 :
(key == 11'b01101011100) ? 46'b1001000001001111110000010010000010011111100000 :
(key == 11'b01101011101) ? 46'b1001000000110100100101010010000001101001001010 :
(key == 11'b01101011110) ? 46'b1001000000011001011011010010000000110010110110 :
(key == 11'b01101011111) ? 46'b1000111111111110010010010001111111111100100100 :
(key == 11'b01101100000) ? 46'b1000111111100011001011110001111111000110010111 :
(key == 11'b01101100001) ? 46'b1000111111001000000101110001111110010000001011 :
(key == 11'b01101100010) ? 46'b1000111110101101000001010001111101011010000010 :
(key == 11'b01101100011) ? 46'b1000111110010001111100110001111100100011111001 :
(key == 11'b01101100100) ? 46'b1000111101110110111100010001111011101101111000 :
(key == 11'b01101100101) ? 46'b1000111101011011111011010001111010110111110110 :
(key == 11'b01101100110) ? 46'b1000111101000000111100110001111010000001111001 :
(key == 11'b01101100111) ? 46'b1000111100100101111111010001111001001011111110 :
(key == 11'b01101101000) ? 46'b1000111100001011000010010001111000010110000100 :
(key == 11'b01101101001) ? 46'b1000111011110000001000010001110111100000010000 :
(key == 11'b01101101010) ? 46'b1000111011010101001110010001110110101010011100 :
(key == 11'b01101101011) ? 46'b1000111010111010010100110001110101110100101001 :
(key == 11'b01101101100) ? 46'b1000111010011111011101110001110100111110111011 :
(key == 11'b01101101101) ? 46'b1000111010000100101001010001110100001001010010 :
(key == 11'b01101101110) ? 46'b1000111001101001110101010001110011010011101010 :
(key == 11'b01101101111) ? 46'b1000111001001111000010010001110010011110000100 :
(key == 11'b01101110000) ? 46'b1000111000110100010000010001110001101000100000 :
(key == 11'b01101110001) ? 46'b1000111000011001100000010001110000110011000000 :
(key == 11'b01101110010) ? 46'b1000110111111110110001010001101111111101100010 :
(key == 11'b01101110011) ? 46'b1000110111100100000011110001101111001000000111 :
(key == 11'b01101110100) ? 46'b1000110111001001011000010001101110010010110000 :
(key == 11'b01101110101) ? 46'b1000110110101110101101010001101101011101011010 :
(key == 11'b01101110110) ? 46'b1000110110010100000011010001101100101000000110 :
(key == 11'b01101110111) ? 46'b1000110101111001011011010001101011110010110110 :
(key == 11'b01101111000) ? 46'b1000110101011110110101010001101010111101101010 :
(key == 11'b01101111001) ? 46'b1000110101000100001111010001101010001000011110 :
(key == 11'b01101111010) ? 46'b1000110100101001101011010001101001010011010110 :
(key == 11'b01101111011) ? 46'b1000110100001111001000010001101000011110010000 :
(key == 11'b01101111100) ? 46'b1000110011110100100111010001100111101001001110 :
(key == 11'b01101111101) ? 46'b1000110011011010000111010001100110110100001110 :
(key == 11'b01101111110) ? 46'b1000110010111111101000010001100101111111010000 :
(key == 11'b01101111111) ? 46'b1000110010100101001010010001100101001010010100 :
(key == 11'b01110000000) ? 46'b1000110010001010101110110001100100010101011101 :
(key == 11'b01110000001) ? 46'b1000110001110000010011010001100011100000100110 :
(key == 11'b01110000010) ? 46'b1000110001010101111001110001100010101011110011 :
(key == 11'b01110000011) ? 46'b1000110000111011100001010001100001110111000010 :
(key == 11'b01110000100) ? 46'b1000110000100001001011010001100001000010010110 :
(key == 11'b01110000101) ? 46'b1000110000000110110110010001100000001101101100 :
(key == 11'b01110000110) ? 46'b1000101111101100100001110001011111011001000011 :
(key == 11'b01110000111) ? 46'b1000101111010010001110010001011110100100011100 :
(key == 11'b01110001000) ? 46'b1000101110110111111100010001011101101111111000 :
(key == 11'b01110001001) ? 46'b1000101110011101101011110001011100111011010111 :
(key == 11'b01110001010) ? 46'b1000101110000011011101010001011100000110111010 :
(key == 11'b01110001011) ? 46'b1000101101101001001111010001011011010010011110 :
(key == 11'b01110001100) ? 46'b1000101101001111000011010001011010011110000110 :
(key == 11'b01110001101) ? 46'b1000101100110100111000010001011001101001110000 :
(key == 11'b01110001110) ? 46'b1000101100011010101110010001011000110101011100 :
(key == 11'b01110001111) ? 46'b1000101100000000100110010001011000000001001100 :
(key == 11'b01110010000) ? 46'b1000101011100110011110010001010111001100111100 :
(key == 11'b01110010001) ? 46'b1000101011001100011000110001010110011000110001 :
(key == 11'b01110010010) ? 46'b1000101010110010010100110001010101100100101001 :
(key == 11'b01110010011) ? 46'b1000101010011000010001010001010100110000100010 :
(key == 11'b01110010100) ? 46'b1000101001111110001111010001010011111100011110 :
(key == 11'b01110010101) ? 46'b1000101001100100001110010001010011001000011100 :
(key == 11'b01110010110) ? 46'b1000101001001010001110010001010010010100011100 :
(key == 11'b01110010111) ? 46'b1000101000110000010000010001010001100000100000 :
(key == 11'b01110011000) ? 46'b1000101000010110010011010001010000101100100110 :
(key == 11'b01110011001) ? 46'b1000100111111100010111010001001111111000101110 :
(key == 11'b01110011010) ? 46'b1000100111100010011110010001001111000100111100 :
(key == 11'b01110011011) ? 46'b1000100111001000100100010001001110010001001000 :
(key == 11'b01110011100) ? 46'b1000100110101110101100010001001101011101011000 :
(key == 11'b01110011101) ? 46'b1000100110010100110110110001001100101001101101 :
(key == 11'b01110011110) ? 46'b1000100101111011000001010001001011110110000010 :
(key == 11'b01110011111) ? 46'b1000100101100001001101010001001011000010011010 :
(key == 11'b01110100000) ? 46'b1000100101000111011010110001001010001110110101 :
(key == 11'b01110100001) ? 46'b1000100100101101101000110001001001011011010001 :
(key == 11'b01110100010) ? 46'b1000100100010011111000010001001000100111110000 :
(key == 11'b01110100011) ? 46'b1000100011111010001010010001000111110100010100 :
(key == 11'b01110100100) ? 46'b1000100011100000011100010001000111000000111000 :
(key == 11'b01110100101) ? 46'b1000100011000110101111110001000110001101011111 :
(key == 11'b01110100110) ? 46'b1000100010101101000100010001000101011010001000 :
(key == 11'b01110100111) ? 46'b1000100010010011011010010001000100100110110100 :
(key == 11'b01110101000) ? 46'b1000100001111001110001110001000011110011100011 :
(key == 11'b01110101001) ? 46'b1000100001100000001011010001000011000000010110 :
(key == 11'b01110101010) ? 46'b1000100001000110100101010001000010001101001010 :
(key == 11'b01110101011) ? 46'b1000100000101101000000010001000001011010000000 :
(key == 11'b01110101100) ? 46'b1000100000010011011100110001000000100110111001 :
(key == 11'b01110101101) ? 46'b1000011111111001111010010000111111110011110100 :
(key == 11'b01110101110) ? 46'b1000011111100000011001010000111111000000110010 :
(key == 11'b01110101111) ? 46'b1000011111000110111001010000111110001101110010 :
(key == 11'b01110110000) ? 46'b1000011110101101011010010000111101011010110100 :
(key == 11'b01110110001) ? 46'b1000011110010011111101010000111100100111111010 :
(key == 11'b01110110010) ? 46'b1000011101111010100001010000111011110101000010 :
(key == 11'b01110110011) ? 46'b1000011101100001000110010000111011000010001100 :
(key == 11'b01110110100) ? 46'b1000011101000111101100010000111010001111011000 :
(key == 11'b01110110101) ? 46'b1000011100101110010100010000111001011100101000 :
(key == 11'b01110110110) ? 46'b1000011100010100111101110000111000101001111011 :
(key == 11'b01110110111) ? 46'b1000011011111011100111010000110111110111001110 :
(key == 11'b01110111000) ? 46'b1000011011100010010010110000110111000100100101 :
(key == 11'b01110111001) ? 46'b1000011011001000111111010000110110010001111110 :
(key == 11'b01110111010) ? 46'b1000011010101111101101010000110101011111011010 :
(key == 11'b01110111011) ? 46'b1000011010010110011011010000110100101100110110 :
(key == 11'b01110111100) ? 46'b1000011001111101001011110000110011111010010111 :
(key == 11'b01110111101) ? 46'b1000011001100011111101110000110011000111111011 :
(key == 11'b01110111110) ? 46'b1000011001001010110000010000110010010101100000 :
(key == 11'b01110111111) ? 46'b1000011000110001100100010000110001100011001000 :
(key == 11'b01111000000) ? 46'b1000011000011000011001010000110000110000110010 :
(key == 11'b01111000001) ? 46'b1000010111111111001110110000101111111110011101 :
(key == 11'b01111000010) ? 46'b1000010111100110000110110000101111001100001101 :
(key == 11'b01111000011) ? 46'b1000010111001100111110110000101110011001111101 :
(key == 11'b01111000100) ? 46'b1000010110110011111001010000101101100111110010 :
(key == 11'b01111000101) ? 46'b1000010110011010110100110000101100110101101001 :
(key == 11'b01111000110) ? 46'b1000010110000001110000010000101100000011100000 :
(key == 11'b01111000111) ? 46'b1000010101101000101101110000101011010001011011 :
(key == 11'b01111001000) ? 46'b1000010101001111101101010000101010011111011010 :
(key == 11'b01111001001) ? 46'b1000010100110110101100110000101001101101011001 :
(key == 11'b01111001010) ? 46'b1000010100011101101101110000101000111011011011 :
(key == 11'b01111001011) ? 46'b1000010100000100110000010000101000001001100000 :
(key == 11'b01111001100) ? 46'b1000010011101011110011010000100111010111100110 :
(key == 11'b01111001101) ? 46'b1000010011010010111000010000100110100101110000 :
(key == 11'b01111001110) ? 46'b1000010010111001111111010000100101110011111110 :
(key == 11'b01111001111) ? 46'b1000010010100001000110010000100101000010001100 :
(key == 11'b01111010000) ? 46'b1000010010001000001110010000100100010000011100 :
(key == 11'b01111010001) ? 46'b1000010001101111011000110000100011011110110001 :
(key == 11'b01111010010) ? 46'b1000010001010110100010110000100010101101000101 :
(key == 11'b01111010011) ? 46'b1000010000111101101111010000100001111011011110 :
(key == 11'b01111010100) ? 46'b1000010000100100111100010000100001001001111000 :
(key == 11'b01111010101) ? 46'b1000010000001100001010010000100000011000010100 :
(key == 11'b01111010110) ? 46'b1000001111110011011001110000011111100110110011 :
(key == 11'b01111010111) ? 46'b1000001111011010101001110000011110110101010011 :
(key == 11'b01111011000) ? 46'b1000001111000001111100110000011110000011111001 :
(key == 11'b01111011001) ? 46'b1000001110101001001111110000011101010010011111 :
(key == 11'b01111011010) ? 46'b1000001110010000100011010000011100100001000110 :
(key == 11'b01111011011) ? 46'b1000001101110111111000110000011011101111110001 :
(key == 11'b01111011100) ? 46'b1000001101011111001111010000011010111110011110 :
(key == 11'b01111011101) ? 46'b1000001101000110100111010000011010001101001110 :
(key == 11'b01111011110) ? 46'b1000001100101110000000010000011001011100000000 :
(key == 11'b01111011111) ? 46'b1000001100010101011010010000011000101010110100 :
(key == 11'b01111100000) ? 46'b1000001011111100110110010000010111111001101100 :
(key == 11'b01111100001) ? 46'b1000001011100100010010010000010111001000100100 :
(key == 11'b01111100010) ? 46'b1000001011001011110000010000010110010111100000 :
(key == 11'b01111100011) ? 46'b1000001010110011001111010000010101100110011110 :
(key == 11'b01111100100) ? 46'b1000001010011010101110110000010100110101011101 :
(key == 11'b01111100101) ? 46'b1000001010000010010000010000010100000100100000 :
(key == 11'b01111100110) ? 46'b1000001001101001110010010000010011010011100100 :
(key == 11'b01111100111) ? 46'b1000001001010001010101010000010010100010101010 :
(key == 11'b01111101000) ? 46'b1000001000111000111001110000010001110001110011 :
(key == 11'b01111101001) ? 46'b1000001000100000011111010000010001000000111110 :
(key == 11'b01111101010) ? 46'b1000001000001000000110010000010000010000001100 :
(key == 11'b01111101011) ? 46'b1000000111101111101110110000001111011111011101 :
(key == 11'b01111101100) ? 46'b1000000111010111011000010000001110101110110000 :
(key == 11'b01111101101) ? 46'b1000000110111111000010010000001101111110000100 :
(key == 11'b01111101110) ? 46'b1000000110100110101101010000001101001101011010 :
(key == 11'b01111101111) ? 46'b1000000110001110011010110000001100011100110101 :
(key == 11'b01111110000) ? 46'b1000000101110110001000110000001011101100010001 :
(key == 11'b01111110001) ? 46'b1000000101011101110111010000001010111011101110 :
(key == 11'b01111110010) ? 46'b1000000101000101100111110000001010001011001111 :
(key == 11'b01111110011) ? 46'b1000000100101101011000110000001001011010110001 :
(key == 11'b01111110100) ? 46'b1000000100010101001011010000001000101010010110 :
(key == 11'b01111110101) ? 46'b1000000011111100111110010000000111111001111100 :
(key == 11'b01111110110) ? 46'b1000000011100100110011010000000111001001100110 :
(key == 11'b01111110111) ? 46'b1000000011001100101001010000000110011001010010 :
(key == 11'b01111111000) ? 46'b1000000010110100100000010000000101101001000000 :
(key == 11'b01111111001) ? 46'b1000000010011100011000010000000100111000110000 :
(key == 11'b01111111010) ? 46'b1000000010000100010001010000000100001000100010 :
(key == 11'b01111111011) ? 46'b1000000001101100001011010000000011011000010110 :
(key == 11'b01111111100) ? 46'b1000000001010100000111110000000010101000001111 :
(key == 11'b01111111101) ? 46'b1000000000111100000100010000000001111000001000 :
(key == 11'b01111111110) ? 46'b1000000000100100000001110000000001001000000011 :
(key == 11'b01111111111) ? 46'b1000000000001100000000010000000000011000000000 :
(key == 11'b10000000000) ? 46'b0000111101110110011110000001111011101100111100 :
(key == 11'b10000000001) ? 46'b0000111101010100100101000001111010101001001010 :
(key == 11'b10000000010) ? 46'b0000111100110010101111000001111001100101011110 :
(key == 11'b10000000011) ? 46'b0000111100010000111100000001111000100001111000 :
(key == 11'b10000000100) ? 46'b0000111011101111001100100001110111011110011001 :
(key == 11'b10000000101) ? 46'b0000111011001101100000100001110110011011000001 :
(key == 11'b10000000110) ? 46'b0000111010101011110111000001110101010111101110 :
(key == 11'b10000000111) ? 46'b0000111010001010010001000001110100010100100010 :
(key == 11'b10000001000) ? 46'b0000111001101000101110000001110011010001011100 :
(key == 11'b10000001001) ? 46'b0000111001000111001110000001110010001110011100 :
(key == 11'b10000001010) ? 46'b0000111000100101110001000001110001001011100010 :
(key == 11'b10000001011) ? 46'b0000111000000100010111100001110000001000101111 :
(key == 11'b10000001100) ? 46'b0000110111100011000000100001101111000110000001 :
(key == 11'b10000001101) ? 46'b0000110111000001101101000001101110000011011010 :
(key == 11'b10000001110) ? 46'b0000110110100000011100100001101101000000111001 :
(key == 11'b10000001111) ? 46'b0000110101111111001111100001101011111110011111 :
(key == 11'b10000010000) ? 46'b0000110101011110000101000001101010111100001010 :
(key == 11'b10000010001) ? 46'b0000110100111100111110000001101001111001111100 :
(key == 11'b10000010010) ? 46'b0000110100011011111010000001101000110111110100 :
(key == 11'b10000010011) ? 46'b0000110011111010111000100001100111110101110001 :
(key == 11'b10000010100) ? 46'b0000110011011001111011000001100110110011110110 :
(key == 11'b10000010101) ? 46'b0000110010111000111111000001100101110001111110 :
(key == 11'b10000010110) ? 46'b0000110010011000000111100001100100110000001111 :
(key == 11'b10000010111) ? 46'b0000110001110111010010000001100011101110100100 :
(key == 11'b10000011000) ? 46'b0000110001010110100000000001100010101101000000 :
(key == 11'b10000011001) ? 46'b0000110000110101110001100001100001101011100011 :
(key == 11'b10000011010) ? 46'b0000110000010101000101000001100000101010001010 :
(key == 11'b10000011011) ? 46'b0000101111110100011100000001011111101000111000 :
(key == 11'b10000011100) ? 46'b0000101111010011110110000001011110100111101100 :
(key == 11'b10000011101) ? 46'b0000101110110011010011000001011101100110100110 :
(key == 11'b10000011110) ? 46'b0000101110010010110010100001011100100101100101 :
(key == 11'b10000011111) ? 46'b0000101101110010010110000001011011100100101100 :
(key == 11'b10000100000) ? 46'b0000101101010001111011000001011010100011110110 :
(key == 11'b10000100001) ? 46'b0000101100110001100100000001011001100011001000 :
(key == 11'b10000100010) ? 46'b0000101100010001001111100001011000100010011111 :
(key == 11'b10000100011) ? 46'b0000101011110000111110000001010111100001111100 :
(key == 11'b10000100100) ? 46'b0000101011010000101111100001010110100001011111 :
(key == 11'b10000100101) ? 46'b0000101010110000100100000001010101100001001000 :
(key == 11'b10000100110) ? 46'b0000101010010000011011000001010100100000110110 :
(key == 11'b10000100111) ? 46'b0000101001110000010110000001010011100000101100 :
(key == 11'b10000101000) ? 46'b0000101001010000010010100001010010100000100101 :
(key == 11'b10000101001) ? 46'b0000101000110000010011000001010001100000100110 :
(key == 11'b10000101010) ? 46'b0000101000010000010110000001010000100000101100 :
(key == 11'b10000101011) ? 46'b0000100111110000011011100001001111100000110111 :
(key == 11'b10000101100) ? 46'b0000100111010000100011100001001110100001000111 :
(key == 11'b10000101101) ? 46'b0000100110110000101111000001001101100001011110 :
(key == 11'b10000101110) ? 46'b0000100110010000111101000001001100100001111010 :
(key == 11'b10000101111) ? 46'b0000100101110001001111000001001011100010011110 :
(key == 11'b10000110000) ? 46'b0000100101010001100011000001001010100011000110 :
(key == 11'b10000110001) ? 46'b0000100100110001111001100001001001100011110011 :
(key == 11'b10000110010) ? 46'b0000100100010010010011000001001000100100100110 :
(key == 11'b10000110011) ? 46'b0000100011110010110000000001000111100101100000 :
(key == 11'b10000110100) ? 46'b0000100011010011001111100001000110100110011111 :
(key == 11'b10000110101) ? 46'b0000100010110011110001100001000101100111100011 :
(key == 11'b10000110110) ? 46'b0000100010010100010110000001000100101000101100 :
(key == 11'b10000110111) ? 46'b0000100001110100111110000001000011101001111100 :
(key == 11'b10000111000) ? 46'b0000100001010101101000100001000010101011010001 :
(key == 11'b10000111001) ? 46'b0000100000110110010110000001000001101100101100 :
(key == 11'b10000111010) ? 46'b0000100000010111000101100001000000101110001011 :
(key == 11'b10000111011) ? 46'b0000011111110111111000100000111111101111110001 :
(key == 11'b10000111100) ? 46'b0000011111011000101110000000111110110001011100 :
(key == 11'b10000111101) ? 46'b0000011110111001100111000000111101110011001110 :
(key == 11'b10000111110) ? 46'b0000011110011010100010000000111100110101000100 :
(key == 11'b10000111111) ? 46'b0000011101111011100000000000111011110111000000 :
(key == 11'b10001000000) ? 46'b0000011101011100100000100000111010111001000001 :
(key == 11'b10001000001) ? 46'b0000011100111101100011000000111001111011000110 :
(key == 11'b10001000010) ? 46'b0000011100011110101001100000111000111101010011 :
(key == 11'b10001000011) ? 46'b0000011011111111110010100000110111111111100101 :
(key == 11'b10001000100) ? 46'b0000011011100000111101100000110111000001111011 :
(key == 11'b10001000101) ? 46'b0000011011000010001100000000110110000100011000 :
(key == 11'b10001000110) ? 46'b0000011010100011011101000000110101000110111010 :
(key == 11'b10001000111) ? 46'b0000011010000100110000100000110100001001100001 :
(key == 11'b10001001000) ? 46'b0000011001100110000111000000110011001100001110 :
(key == 11'b10001001001) ? 46'b0000011001000111011111100000110010001110111111 :
(key == 11'b10001001010) ? 46'b0000011000101000111011100000110001010001110111 :
(key == 11'b10001001011) ? 46'b0000011000001010011010000000110000010100110100 :
(key == 11'b10001001100) ? 46'b0000010111101011111010100000101111010111110101 :
(key == 11'b10001001101) ? 46'b0000010111001101011110000000101110011010111100 :
(key == 11'b10001001110) ? 46'b0000010110101111000100000000101101011110001000 :
(key == 11'b10001001111) ? 46'b0000010110010000101101100000101100100001011011 :
(key == 11'b10001010000) ? 46'b0000010101110010011001000000101011100100110010 :
(key == 11'b10001010001) ? 46'b0000010101010100000111000000101010101000001110 :
(key == 11'b10001010010) ? 46'b0000010100110101111000000000101001101011110000 :
(key == 11'b10001010011) ? 46'b0000010100010111101011100000101000101111010111 :
(key == 11'b10001010100) ? 46'b0000010011111001100001000000100111110011000010 :
(key == 11'b10001010101) ? 46'b0000010011011011011010000000100110110110110100 :
(key == 11'b10001010110) ? 46'b0000010010111101010101000000100101111010101010 :
(key == 11'b10001010111) ? 46'b0000010010011111010011000000100100111110100110 :
(key == 11'b10001011000) ? 46'b0000010010000001010100000000100100000010101000 :
(key == 11'b10001011001) ? 46'b0000010001100011010111000000100011000110101110 :
(key == 11'b10001011010) ? 46'b0000010001000101011100000000100010001010111000 :
(key == 11'b10001011011) ? 46'b0000010000100111100100000000100001001111001000 :
(key == 11'b10001011100) ? 46'b0000010000001001101111000000100000010011011110 :
(key == 11'b10001011101) ? 46'b0000001111101011111100000000011111010111111000 :
(key == 11'b10001011110) ? 46'b0000001111001110001100000000011110011100011000 :
(key == 11'b10001011111) ? 46'b0000001110110000011111000000011101100000111110 :
(key == 11'b10001100000) ? 46'b0000001110010010110100000000011100100101101000 :
(key == 11'b10001100001) ? 46'b0000001101110101001011100000011011101010010111 :
(key == 11'b10001100010) ? 46'b0000001101010111100101000000011010101111001010 :
(key == 11'b10001100011) ? 46'b0000001100111010000010000000011001110100000100 :
(key == 11'b10001100100) ? 46'b0000001100011100100001000000011000111001000010 :
(key == 11'b10001100101) ? 46'b0000001011111111000010100000010111111110000101 :
(key == 11'b10001100110) ? 46'b0000001011100001100111000000010111000011001110 :
(key == 11'b10001100111) ? 46'b0000001011000100001101000000010110001000011010 :
(key == 11'b10001101000) ? 46'b0000001010100110110110100000010101001101101101 :
(key == 11'b10001101001) ? 46'b0000001010001001100010100000010100010011000101 :
(key == 11'b10001101010) ? 46'b0000001001101100010000100000010011011000100001 :
(key == 11'b10001101011) ? 46'b0000001001001111000001000000010010011110000010 :
(key == 11'b10001101100) ? 46'b0000001000110001110100000000010001100011101000 :
(key == 11'b10001101101) ? 46'b0000001000010100101001100000010000101001010011 :
(key == 11'b10001101110) ? 46'b0000000111110111100010000000001111101111000100 :
(key == 11'b10001101111) ? 46'b0000000111011010011100000000001110110100111000 :
(key == 11'b10001110000) ? 46'b0000000110111101011001000000001101111010110010 :
(key == 11'b10001110001) ? 46'b0000000110100000011000100000001101000000110001 :
(key == 11'b10001110010) ? 46'b0000000110000011011010100000001100000110110101 :
(key == 11'b10001110011) ? 46'b0000000101100110011111000000001011001100111110 :
(key == 11'b10001110100) ? 46'b0000000101001001100101100000001010010011001011 :
(key == 11'b10001110101) ? 46'b0000000100101100101110100000001001011001011101 :
(key == 11'b10001110110) ? 46'b0000000100001111111010000000001000011111110100 :
(key == 11'b10001110111) ? 46'b0000000011110011001000000000000111100110010000 :
(key == 11'b10001111000) ? 46'b0000000011010110011000100000000110101100110001 :
(key == 11'b10001111001) ? 46'b0000000010111001101011100000000101110011010111 :
(key == 11'b10001111010) ? 46'b0000000010011101000000100000000100111010000001 :
(key == 11'b10001111011) ? 46'b0000000010000000011000000000000100000000110000 :
(key == 11'b10001111100) ? 46'b0000000001100011110010100000000011000111100101 :
(key == 11'b10001111101) ? 46'b0000000001000111001111000000000010001110011110 :
(key == 11'b10001111110) ? 46'b0000000000101010101101100000000001010101011011 :
(key == 11'b10001111111) ? 46'b0000000000001110001111000000000000011100011110 :
(key == 11'b10010000000) ? 46'b1111111111100011100101011111111111000111001010 :
(key == 11'b10010000001) ? 46'b1111111110101010110000011111111101010101100000 :
(key == 11'b10010000010) ? 46'b1111111101110010000001011111111011100100000010 :
(key == 11'b10010000011) ? 46'b1111111100111001010111011111111001110010101110 :
(key == 11'b10010000100) ? 46'b1111111100000000110000111111111000000001100001 :
(key == 11'b10010000101) ? 46'b1111111011001000001111011111110110010000011110 :
(key == 11'b10010000110) ? 46'b1111111010001111110010111111110100011111100101 :
(key == 11'b10010000111) ? 46'b1111111001010111011011011111110010101110110110 :
(key == 11'b10010001000) ? 46'b1111111000011111001000011111110000111110010000 :
(key == 11'b10010001001) ? 46'b1111110111100110111001111111101111001101110011 :
(key == 11'b10010001010) ? 46'b1111110110101110101111011111101101011101011110 :
(key == 11'b10010001011) ? 46'b1111110101110110101001011111101011101101010010 :
(key == 11'b10010001100) ? 46'b1111110100111110101001011111101001111101010010 :
(key == 11'b10010001101) ? 46'b1111110100000110101100111111101000001101011001 :
(key == 11'b10010001110) ? 46'b1111110011001110110100111111100110011101101001 :
(key == 11'b10010001111) ? 46'b1111110010010111000010011111100100101110000100 :
(key == 11'b10010010000) ? 46'b1111110001011111010011111111100010111110100111 :
(key == 11'b10010010001) ? 46'b1111110000100111101010011111100001001111010100 :
(key == 11'b10010010010) ? 46'b1111101111110000000100111111011111100000001001 :
(key == 11'b10010010011) ? 46'b1111101110111000100100011111011101110001001000 :
(key == 11'b10010010100) ? 46'b1111101110000001000111111111011100000010001111 :
(key == 11'b10010010101) ? 46'b1111101101001001110000111111011010010011100001 :
(key == 11'b10010010110) ? 46'b1111101100010010011101011111011000100100111010 :
(key == 11'b10010010111) ? 46'b1111101011011011001110111111010110110110011101 :
(key == 11'b10010011000) ? 46'b1111101010100100000101011111010101001000001010 :
(key == 11'b10010011001) ? 46'b1111101001101101000000011111010011011010000000 :
(key == 11'b10010011010) ? 46'b1111101000110101111111011111010001101011111110 :
(key == 11'b10010011011) ? 46'b1111100111111111000010011111001111111110000100 :
(key == 11'b10010011100) ? 46'b1111100111001000001010011111001110010000010100 :
(key == 11'b10010011101) ? 46'b1111100110010001010110011111001100100010101100 :
(key == 11'b10010011110) ? 46'b1111100101011010100111111111001010110101001111 :
(key == 11'b10010011111) ? 46'b1111100100100011111100011111001001000111111000 :
(key == 11'b10010100000) ? 46'b1111100011101101010110111111000111011010101101 :
(key == 11'b10010100001) ? 46'b1111100010110110110100011111000101101101101000 :
(key == 11'b10010100010) ? 46'b1111100010000000010111011111000100000000101110 :
(key == 11'b10010100011) ? 46'b1111100001001001111110011111000010010011111100 :
(key == 11'b10010100100) ? 46'b1111100000010011101001011111000000100111010010 :
(key == 11'b10010100101) ? 46'b1111011111011101011000111110111110111010110001 :
(key == 11'b10010100110) ? 46'b1111011110100111001100111110111101001110011001 :
(key == 11'b10010100111) ? 46'b1111011101110001000101011110111011100010001010 :
(key == 11'b10010101000) ? 46'b1111011100111011000010011110111001110110000100 :
(key == 11'b10010101001) ? 46'b1111011100000101000011111110111000001010000111 :
(key == 11'b10010101010) ? 46'b1111011011001111001001011110110110011110010010 :
(key == 11'b10010101011) ? 46'b1111011010011001010010111110110100110010100101 :
(key == 11'b10010101100) ? 46'b1111011001100011100001011110110011000111000010 :
(key == 11'b10010101101) ? 46'b1111011000101101110011111110110001011011100111 :
(key == 11'b10010101110) ? 46'b1111010111111000001010011110101111110000010100 :
(key == 11'b10010101111) ? 46'b1111010111000010100101011110101110000101001010 :
(key == 11'b10010110000) ? 46'b1111010110001101000100111110101100011010001001 :
(key == 11'b10010110001) ? 46'b1111010101010111101000111110101010101111010001 :
(key == 11'b10010110010) ? 46'b1111010100100010001111111110101001000100011111 :
(key == 11'b10010110011) ? 46'b1111010011101100111100011110100111011001111000 :
(key == 11'b10010110100) ? 46'b1111010010110111101100111110100101101111011001 :
(key == 11'b10010110101) ? 46'b1111010010000010100001011110100100000101000010 :
(key == 11'b10010110110) ? 46'b1111010001001101011010011110100010011010110100 :
(key == 11'b10010110111) ? 46'b1111010000011000010111111110100000110000101111 :
(key == 11'b10010111000) ? 46'b1111001111100011011000011110011111000110110000 :
(key == 11'b10010111001) ? 46'b1111001110101110011110011110011101011100111100 :
(key == 11'b10010111010) ? 46'b1111001101111001101000011110011011110011010000 :
(key == 11'b10010111011) ? 46'b1111001101000100110110011110011010001001101100 :
(key == 11'b10010111100) ? 46'b1111001100010000001000011110011000100000010000 :
(key == 11'b10010111101) ? 46'b1111001011011011011110011110010110110110111100 :
(key == 11'b10010111110) ? 46'b1111001010100110111001011110010101001101110010 :
(key == 11'b10010111111) ? 46'b1111001001110010010111011110010011100100101110 :
(key == 11'b10011000000) ? 46'b1111001000111101111001111110010001111011110011 :
(key == 11'b10011000001) ? 46'b1111001000001001100001011110010000010011000010 :
(key == 11'b10011000010) ? 46'b1111000111010101001011111110001110101010010111 :
(key == 11'b10011000011) ? 46'b1111000110100000111010111110001101000001110101 :
(key == 11'b10011000100) ? 46'b1111000101101100101110011110001011011001011100 :
(key == 11'b10011000101) ? 46'b1111000100111000100110011110001001110001001100 :
(key == 11'b10011000110) ? 46'b1111000100000100100001011110001000001001000010 :
(key == 11'b10011000111) ? 46'b1111000011010000100000111110000110100001000001 :
(key == 11'b10011001000) ? 46'b1111000010011100100100011110000100111001001000 :
(key == 11'b10011001001) ? 46'b1111000001101000101011111110000011010001010111 :
(key == 11'b10011001010) ? 46'b1111000000110100110111011110000001101001101110 :
(key == 11'b10011001011) ? 46'b1111000000000001000111011110000000000010001110 :
(key == 11'b10011001100) ? 46'b1110111111001101011011011101111110011010110110 :
(key == 11'b10011001101) ? 46'b1110111110011001110011011101111100110011100110 :
(key == 11'b10011001110) ? 46'b1110111101100110001111011101111011001100011110 :
(key == 11'b10011001111) ? 46'b1110111100110010101111011101111001100101011110 :
(key == 11'b10011010000) ? 46'b1110111011111111010011011101110111111110100110 :
(key == 11'b10011010001) ? 46'b1110111011001011111010011101110110010111110100 :
(key == 11'b10011010010) ? 46'b1110111010011000100110011101110100110001001100 :
(key == 11'b10011010011) ? 46'b1110111001100101010111011101110011001010101110 :
(key == 11'b10011010100) ? 46'b1110111000110010001010011101110001100100010100 :
(key == 11'b10011010101) ? 46'b1110110111111111000010011101101111111110000100 :
(key == 11'b10011010110) ? 46'b1110110111001011111101111101101110010111111011 :
(key == 11'b10011010111) ? 46'b1110110110011000111101111101101100110001111011 :
(key == 11'b10011011000) ? 46'b1110110101100110000001011101101011001100000010 :
(key == 11'b10011011001) ? 46'b1110110100110011001001011101101001100110010010 :
(key == 11'b10011011010) ? 46'b1110110100000000010100011101101000000000101000 :
(key == 11'b10011011011) ? 46'b1110110011001101100100111101100110011011001001 :
(key == 11'b10011011100) ? 46'b1110110010011010111000011101100100110101110000 :
(key == 11'b10011011101) ? 46'b1110110001101000001110111101100011010000011101 :
(key == 11'b10011011110) ? 46'b1110110000110101101001111101100001101011010011 :
(key == 11'b10011011111) ? 46'b1110110000000011001001011101100000000110010010 :
(key == 11'b10011100000) ? 46'b1110101111010000101101011101011110100001011010 :
(key == 11'b10011100001) ? 46'b1110101110011110010011011101011100111100100110 :
(key == 11'b10011100010) ? 46'b1110101101101011111110011101011011010111111100 :
(key == 11'b10011100011) ? 46'b1110101100111001101100111101011001110011011001 :
(key == 11'b10011100100) ? 46'b1110101100000111011111111101011000001110111111 :
(key == 11'b10011100101) ? 46'b1110101011010101010101111101010110101010101011 :
(key == 11'b10011100110) ? 46'b1110101010100011010000011101010101000110100000 :
(key == 11'b10011100111) ? 46'b1110101001110001001101111101010011100010011011 :
(key == 11'b10011101000) ? 46'b1110101000111111001111111101010001111110011111 :
(key == 11'b10011101001) ? 46'b1110101000001101010101011101010000011010101010 :
(key == 11'b10011101010) ? 46'b1110100111011011011111011101001110110110111110 :
(key == 11'b10011101011) ? 46'b1110100110101001101100011101001101010011011000 :
(key == 11'b10011101100) ? 46'b1110100101110111111101011101001011101111111010 :
(key == 11'b10011101101) ? 46'b1110100101000110010010011101001010001100100100 :
(key == 11'b10011101110) ? 46'b1110100100010100101011011101001000101001010110 :
(key == 11'b10011101111) ? 46'b1110100011100011000110111101000111000110001101 :
(key == 11'b10011110000) ? 46'b1110100010110001100110111101000101100011001101 :
(key == 11'b10011110001) ? 46'b1110100010000000001011011101000100000000010110 :
(key == 11'b10011110010) ? 46'b1110100001001110110010111101000010011101100101 :
(key == 11'b10011110011) ? 46'b1110100000011101011101011101000000111010111010 :
(key == 11'b10011110100) ? 46'b1110011111101100001101011100111111011000011010 :
(key == 11'b10011110101) ? 46'b1110011110111011000000011100111101110110000000 :
(key == 11'b10011110110) ? 46'b1110011110001001110111011100111100010011101110 :
(key == 11'b10011110111) ? 46'b1110011101011000110001011100111010110001100010 :
(key == 11'b10011111000) ? 46'b1110011100100111101110011100111001001111011100 :
(key == 11'b10011111001) ? 46'b1110011011110110110000011100110111101101100000 :
(key == 11'b10011111010) ? 46'b1110011011000101110101111100110110001011101011 :
(key == 11'b10011111011) ? 46'b1110011010010100111111011100110100101001111110 :
(key == 11'b10011111100) ? 46'b1110011001100100001100011100110011001000011000 :
(key == 11'b10011111101) ? 46'b1110011000110011011100011100110001100110111000 :
(key == 11'b10011111110) ? 46'b1110011000000010101111111100110000000101011111 :
(key == 11'b10011111111) ? 46'b1110010111010010000111011100101110100100001110 :
(key == 11'b10100000000) ? 46'b1110010110100001100011011100101101000011000110 :
(key == 11'b10100000001) ? 46'b1110010101110001000010011100101011100010000100 :
(key == 11'b10100000010) ? 46'b1110010101000000100100011100101010000001001000 :
(key == 11'b10100000011) ? 46'b1110010100010000001010111100101000100000010101 :
(key == 11'b10100000100) ? 46'b1110010011011111110100011100100110111111101000 :
(key == 11'b10100000101) ? 46'b1110010010101111100010011100100101011111000100 :
(key == 11'b10100000110) ? 46'b1110010001111111010011011100100011111110100110 :
(key == 11'b10100000111) ? 46'b1110010001001111001000011100100010011110010000 :
(key == 11'b10100001000) ? 46'b1110010000011111000000011100100000111110000000 :
(key == 11'b10100001001) ? 46'b1110001111101110111100111100011111011101111001 :
(key == 11'b10100001010) ? 46'b1110001110111110111011011100011101111101110110 :
(key == 11'b10100001011) ? 46'b1110001110001110111110011100011100011101111100 :
(key == 11'b10100001100) ? 46'b1110001101011111000101111100011010111110001011 :
(key == 11'b10100001101) ? 46'b1110001100101111001110111100011001011110011101 :
(key == 11'b10100001110) ? 46'b1110001011111111011100011100010111111110111000 :
(key == 11'b10100001111) ? 46'b1110001011001111101110011100010110011111011100 :
(key == 11'b10100010000) ? 46'b1110001010100000000010011100010101000000000100 :
(key == 11'b10100010001) ? 46'b1110001001110000011011011100010011100000110110 :
(key == 11'b10100010010) ? 46'b1110001001000000110110011100010010000001101100 :
(key == 11'b10100010011) ? 46'b1110001000010001010101111100010000100010101011 :
(key == 11'b10100010100) ? 46'b1110000111100001111001011100001111000011110010 :
(key == 11'b10100010101) ? 46'b1110000110110010011111011100001101100100111110 :
(key == 11'b10100010110) ? 46'b1110000110000011001001011100001100000110010010 :
(key == 11'b10100010111) ? 46'b1110000101010011110110011100001010100111101100 :
(key == 11'b10100011000) ? 46'b1110000100100100100111111100001001001001001111 :
(key == 11'b10100011001) ? 46'b1110000011110101011011011100000111101010110110 :
(key == 11'b10100011010) ? 46'b1110000011000110010011111100000110001100100111 :
(key == 11'b10100011011) ? 46'b1110000010010111001110011100000100101110011100 :
(key == 11'b10100011100) ? 46'b1110000001101000001101011100000011010000011010 :
(key == 11'b10100011101) ? 46'b1110000000111001001111011100000001110010011110 :
(key == 11'b10100011110) ? 46'b1110000000001010010100011100000000010100101000 :
(key == 11'b10100011111) ? 46'b1101111111011011011101111011111110110110111011 :
(key == 11'b10100100000) ? 46'b1101111110101100101010011011111101011001010100 :
(key == 11'b10100100001) ? 46'b1101111101111101111001111011111011111011110011 :
(key == 11'b10100100010) ? 46'b1101111101001111001101011011111010011110011010 :
(key == 11'b10100100011) ? 46'b1101111100100000100011011011111001000001000110 :
(key == 11'b10100100100) ? 46'b1101111011110001111110011011110111100011111100 :
(key == 11'b10100100101) ? 46'b1101111011000011011011111011110110000110110111 :
(key == 11'b10100100110) ? 46'b1101111010010100111011111011110100101001110111 :
(key == 11'b10100100111) ? 46'b1101111001100110100000011011110011001101000000 :
(key == 11'b10100101000) ? 46'b1101111000111000000111111011110001110000001111 :
(key == 11'b10100101001) ? 46'b1101111000001001110010011011110000010011100100 :
(key == 11'b10100101010) ? 46'b1101110111011011100001011011101110110111000010 :
(key == 11'b10100101011) ? 46'b1101110110101101010010011011101101011010100100 :
(key == 11'b10100101100) ? 46'b1101110101111111001000011011101011111110010000 :
(key == 11'b10100101101) ? 46'b1101110101010001000000011011101010100010000000 :
(key == 11'b10100101110) ? 46'b1101110100100010111100011011101001000101111000 :
(key == 11'b10100101111) ? 46'b1101110011110100111010111011100111101001110101 :
(key == 11'b10100110000) ? 46'b1101110011000110111101011011100110001101111010 :
(key == 11'b10100110001) ? 46'b1101110010011001000010111011100100110010000101 :
(key == 11'b10100110010) ? 46'b1101110001101011001100011011100011010110011000 :
(key == 11'b10100110011) ? 46'b1101110000111101011000011011100001111010110000 :
(key == 11'b10100110100) ? 46'b1101110000001111100111011011100000011111001110 :
(key == 11'b10100110101) ? 46'b1101101111100001111010011011011111000011110100 :
(key == 11'b10100110110) ? 46'b1101101110110100010001011011011101101000100010 :
(key == 11'b10100110111) ? 46'b1101101110000110101010011011011100001101010100 :
(key == 11'b10100111000) ? 46'b1101101101011001000111111011011010110010001111 :
(key == 11'b10100111001) ? 46'b1101101100101011100110111011011001010111001101 :
(key == 11'b10100111010) ? 46'b1101101011111110001010011011010111111100010100 :
(key == 11'b10100111011) ? 46'b1101101011010000110000111011010110100001100001 :
(key == 11'b10100111100) ? 46'b1101101010100011011011011011010101000110110110 :
(key == 11'b10100111101) ? 46'b1101101001110110001000011011010011101100010000 :
(key == 11'b10100111110) ? 46'b1101101001001000110111111011010010010001101111 :
(key == 11'b10100111111) ? 46'b1101101000011011101011111011010000110111010111 :
(key == 11'b10101000000) ? 46'b1101100111101110100010111011001111011101000101 :
(key == 11'b10101000001) ? 46'b1101100111000001011100011011001110000010111000 :
(key == 11'b10101000010) ? 46'b1101100110010100011001111011001100101000110011 :
(key == 11'b10101000011) ? 46'b1101100101100111011001111011001011001110110011 :
(key == 11'b10101000100) ? 46'b1101100100111010011101011011001001110100111010 :
(key == 11'b10101000101) ? 46'b1101100100001101100100011011001000011011001000 :
(key == 11'b10101000110) ? 46'b1101100011100000101110011011000111000001011100 :
(key == 11'b10101000111) ? 46'b1101100010110011111011011011000101100111110110 :
(key == 11'b10101001000) ? 46'b1101100010000111001100011011000100001110011000 :
(key == 11'b10101001001) ? 46'b1101100001011010011110111011000010110100111101 :
(key == 11'b10101001010) ? 46'b1101100000101101110101011011000001011011101010 :
(key == 11'b10101001011) ? 46'b1101100000000001010000011011000000000010100000 :
(key == 11'b10101001100) ? 46'b1101011111010100101100111010111110101001011001 :
(key == 11'b10101001101) ? 46'b1101011110101000001100011010111101010000011000 :
(key == 11'b10101001110) ? 46'b1101011101111011110000011010111011110111100000 :
(key == 11'b10101001111) ? 46'b1101011101001111010111011010111010011110101110 :
(key == 11'b10101010000) ? 46'b1101011100100010111111111010111001000101111111 :
(key == 11'b10101010001) ? 46'b1101011011110110101100111010110111101101011001 :
(key == 11'b10101010010) ? 46'b1101011011001010011100111010110110010100111001 :
(key == 11'b10101010011) ? 46'b1101011010011110001111111010110100111100011111 :
(key == 11'b10101010100) ? 46'b1101011001110010000101111010110011100100001011 :
(key == 11'b10101010101) ? 46'b1101011001000101111110111010110010001011111101 :
(key == 11'b10101010110) ? 46'b1101011000011001111011011010110000110011110110 :
(key == 11'b10101010111) ? 46'b1101010111101101111011011010101111011011110110 :
(key == 11'b10101011000) ? 46'b1101010111000001111101011010101110000011111010 :
(key == 11'b10101011001) ? 46'b1101010110010110000010011010101100101100000100 :
(key == 11'b10101011010) ? 46'b1101010101101010001011111010101011010100010111 :
(key == 11'b10101011011) ? 46'b1101010100111110010110111010101001111100101101 :
(key == 11'b10101011100) ? 46'b1101010100010010100101011010101000100101001010 :
(key == 11'b10101011101) ? 46'b1101010011100110110111011010100111001101101110 :
(key == 11'b10101011110) ? 46'b1101010010111011001100011010100101110110011000 :
(key == 11'b10101011111) ? 46'b1101010010001111100011111010100100011111000111 :
(key == 11'b10101100000) ? 46'b1101010001100011111111011010100011000111111110 :
(key == 11'b10101100001) ? 46'b1101010000111000011100011010100001110000111000 :
(key == 11'b10101100010) ? 46'b1101010000001100111101111010100000011001111011 :
(key == 11'b10101100011) ? 46'b1101001111100001100010011010011111000011000100 :
(key == 11'b10101100100) ? 46'b1101001110110110001001011010011101101100010010 :
(key == 11'b10101100101) ? 46'b1101001110001010110010111010011100010101100101 :
(key == 11'b10101100110) ? 46'b1101001101011111100000011010011010111111000000 :
(key == 11'b10101100111) ? 46'b1101001100110100010000111010011001101000100001 :
(key == 11'b10101101000) ? 46'b1101001100001001000010111010011000010010000101 :
(key == 11'b10101101001) ? 46'b1101001011011101111001011010010110111011110010 :
(key == 11'b10101101010) ? 46'b1101001010110010110010011010010101100101100100 :
(key == 11'b10101101011) ? 46'b1101001010000111101110011010010100001111011100 :
(key == 11'b10101101100) ? 46'b1101001001011100101101011010010010111001011010 :
(key == 11'b10101101101) ? 46'b1101001000110001101111111010010001100011011111 :
(key == 11'b10101101110) ? 46'b1101001000000110110100011010010000001101101000 :
(key == 11'b10101101111) ? 46'b1101000111011011111100011010001110110111111000 :
(key == 11'b10101110000) ? 46'b1101000110110001000111111010001101100010001111 :
(key == 11'b10101110001) ? 46'b1101000110000110010100111010001100001100101001 :
(key == 11'b10101110010) ? 46'b1101000101011011100110011010001010110111001100 :
(key == 11'b10101110011) ? 46'b1101000100110000111001011010001001100001110010 :
(key == 11'b10101110100) ? 46'b1101000100000110010000111010001000001100100001 :
(key == 11'b10101110101) ? 46'b1101000011011011101001111010000110110111010011 :
(key == 11'b10101110110) ? 46'b1101000010110001000101111010000101100010001011 :
(key == 11'b10101110111) ? 46'b1101000010000110100101011010000100001101001010 :
(key == 11'b10101111000) ? 46'b1101000001011100001000011010000010111000010000 :
(key == 11'b10101111001) ? 46'b1101000000110001101101011010000001100011011010 :
(key == 11'b10101111010) ? 46'b1101000000000111010101011010000000001110101010 :
(key == 11'b10101111011) ? 46'b1100111111011101000000011001111110111010000000 :
(key == 11'b10101111100) ? 46'b1100111110110010101110011001111101100101011100 :
(key == 11'b10101111101) ? 46'b1100111110001000011111011001111100010000111110 :
(key == 11'b10101111110) ? 46'b1100111101011110010011011001111010111100100110 :
(key == 11'b10101111111) ? 46'b1100111100110100001001011001111001101000010010 :
(key == 11'b10110000000) ? 46'b1100111100001010000010111001111000010100000101 :
(key == 11'b10110000001) ? 46'b1100111011011111111111111001110110111111111111 :
(key == 11'b10110000010) ? 46'b1100111010110101111110011001110101101011111100 :
(key == 11'b10110000011) ? 46'b1100111010001100000001011001110100011000000010 :
(key == 11'b10110000100) ? 46'b1100111001100010000101111001110011000100001011 :
(key == 11'b10110000101) ? 46'b1100111000111000001101011001110001110000011010 :
(key == 11'b10110000110) ? 46'b1100111000001110010111111001110000011100101111 :
(key == 11'b10110000111) ? 46'b1100110111100100100101011001101111001001001010 :
(key == 11'b10110001000) ? 46'b1100110110111010110101111001101101110101101011 :
(key == 11'b10110001001) ? 46'b1100110110010001001001011001101100100010010010 :
(key == 11'b10110001010) ? 46'b1100110101100111011111011001101011001110111110 :
(key == 11'b10110001011) ? 46'b1100110100111101110111111001101001111011101111 :
(key == 11'b10110001100) ? 46'b1100110100010100010010111001101000101000100101 :
(key == 11'b10110001101) ? 46'b1100110011101010110000111001100111010101100001 :
(key == 11'b10110001110) ? 46'b1100110011000001010010011001100110000010100100 :
(key == 11'b10110001111) ? 46'b1100110010010111110110011001100100101111101100 :
(key == 11'b10110010000) ? 46'b1100110001101110011101011001100011011100111010 :
(key == 11'b10110010001) ? 46'b1100110001000101000110111001100010001010001101 :
(key == 11'b10110010010) ? 46'b1100110000011011110011111001100000110111100111 :
(key == 11'b10110010011) ? 46'b1100101111110010100010011001011111100101000100 :
(key == 11'b10110010100) ? 46'b1100101111001001010100011001011110010010101000 :
(key == 11'b10110010101) ? 46'b1100101110100000001001011001011101000000010010 :
(key == 11'b10110010110) ? 46'b1100101101110110111111111001011011101101111111 :
(key == 11'b10110010111) ? 46'b1100101101001101111010011001011010011011110100 :
(key == 11'b10110011000) ? 46'b1100101100100100110111111001011001001001101111 :
(key == 11'b10110011001) ? 46'b1100101011111011110110111001010111110111101101 :
(key == 11'b10110011010) ? 46'b1100101011010010111001011001010110100101110010 :
(key == 11'b10110011011) ? 46'b1100101010101001111110011001010101010011111100 :
(key == 11'b10110011100) ? 46'b1100101010000001000110011001010100000010001100 :
(key == 11'b10110011101) ? 46'b1100101001011000010001011001010010110000100010 :
(key == 11'b10110011110) ? 46'b1100101000101111011110111001010001011110111101 :
(key == 11'b10110011111) ? 46'b1100101000000110101110011001010000001101011100 :
(key == 11'b10110100000) ? 46'b1100100111011110000001011001001110111100000010 :
(key == 11'b10110100001) ? 46'b1100100110110101010111011001001101101010101110 :
(key == 11'b10110100010) ? 46'b1100100110001100101110111001001100011001011101 :
(key == 11'b10110100011) ? 46'b1100100101100100001010011001001011001000010100 :
(key == 11'b10110100100) ? 46'b1100100100111011100111011001001001110111001110 :
(key == 11'b10110100101) ? 46'b1100100100010011001000011001001000100110010000 :
(key == 11'b10110100110) ? 46'b1100100011101010101011011001000111010101010110 :
(key == 11'b10110100111) ? 46'b1100100011000010010000011001000110000100100000 :
(key == 11'b10110101000) ? 46'b1100100010011001111001011001000100110011110010 :
(key == 11'b10110101001) ? 46'b1100100001110001100011111001000011100011000111 :
(key == 11'b10110101010) ? 46'b1100100001001001010010011001000010010010100100 :
(key == 11'b10110101011) ? 46'b1100100000100001000001111001000001000010000011 :
(key == 11'b10110101100) ? 46'b1100011111111000110101011000111111110001101010 :
(key == 11'b10110101101) ? 46'b1100011111010000101010011000111110100001010100 :
(key == 11'b10110101110) ? 46'b1100011110101000100011011000111101010001000110 :
(key == 11'b10110101111) ? 46'b1100011110000000011110011000111100000000111100 :
(key == 11'b10110110000) ? 46'b1100011101011000011011011000111010110000110110 :
(key == 11'b10110110001) ? 46'b1100011100110000011100011000111001100000111000 :
(key == 11'b10110110010) ? 46'b1100011100001000011110111000111000010000111101 :
(key == 11'b10110110011) ? 46'b1100011011100000100100011000110111000001001000 :
(key == 11'b10110110100) ? 46'b1100011010111000101100111000110101110001011001 :
(key == 11'b10110110101) ? 46'b1100011010010000110110111000110100100001101101 :
(key == 11'b10110110110) ? 46'b1100011001101001000100011000110011010010001000 :
(key == 11'b10110110111) ? 46'b1100011001000001010100011000110010000010101000 :
(key == 11'b10110111000) ? 46'b1100011000011001100110111000110000110011001101 :
(key == 11'b10110111001) ? 46'b1100010111110001111100111000101111100011111001 :
(key == 11'b10110111010) ? 46'b1100010111001010010100011000101110010100101000 :
(key == 11'b10110111011) ? 46'b1100010110100010101110111000101101000101011101 :
(key == 11'b10110111100) ? 46'b1100010101111011001100011000101011110110011000 :
(key == 11'b10110111101) ? 46'b1100010101010011101011011000101010100111010110 :
(key == 11'b10110111110) ? 46'b1100010100101100001101011000101001011000011010 :
(key == 11'b10110111111) ? 46'b1100010100000100110010011000101000001001100100 :
(key == 11'b10111000000) ? 46'b1100010011011101011000111000100110111010110001 :
(key == 11'b10111000001) ? 46'b1100010010110110000011011000100101101100000110 :
(key == 11'b10111000010) ? 46'b1100010010001110101110111000100100011101011101 :
(key == 11'b10111000011) ? 46'b1100010001100111011110011000100011001110111100 :
(key == 11'b10111000100) ? 46'b1100010001000000010000011000100010000000100000 :
(key == 11'b10111000101) ? 46'b1100010000011001000100011000100000110010001000 :
(key == 11'b10111000110) ? 46'b1100001111110001111010011000011111100011110100 :
(key == 11'b10111000111) ? 46'b1100001111001010110011011000011110010101100110 :
(key == 11'b10111001000) ? 46'b1100001110100011101111111000011101000111011111 :
(key == 11'b10111001001) ? 46'b1100001101111100101110011000011011111001011100 :
(key == 11'b10111001010) ? 46'b1100001101010101101110011000011010101011011100 :
(key == 11'b10111001011) ? 46'b1100001100101110110001011000011001011101100010 :
(key == 11'b10111001100) ? 46'b1100001100000111110111011000011000001111101110 :
(key == 11'b10111001101) ? 46'b1100001011100001000000011000010111000010000000 :
(key == 11'b10111001110) ? 46'b1100001010111010001010111000010101110100010101 :
(key == 11'b10111001111) ? 46'b1100001010010011011000011000010100100110110000 :
(key == 11'b10111010000) ? 46'b1100001001101100100111011000010011011001001110 :
(key == 11'b10111010001) ? 46'b1100001001000101111010011000010010001011110100 :
(key == 11'b10111010010) ? 46'b1100001000011111001110011000010000111110011100 :
(key == 11'b10111010011) ? 46'b1100000111111000100110011000001111110001001100 :
(key == 11'b10111010100) ? 46'b1100000111010001111111111000001110100011111111 :
(key == 11'b10111010101) ? 46'b1100000110101011011100011000001101010110111000 :
(key == 11'b10111010110) ? 46'b1100000110000100111011011000001100001001110110 :
(key == 11'b10111010111) ? 46'b1100000101011110011100011000001010111100111000 :
(key == 11'b10111011000) ? 46'b1100000100110111111111011000001001101111111110 :
(key == 11'b10111011001) ? 46'b1100000100010001100110011000001000100011001100 :
(key == 11'b10111011010) ? 46'b1100000011101011001110111000000111010110011101 :
(key == 11'b10111011011) ? 46'b1100000011000100111010011000000110001001110100 :
(key == 11'b10111011100) ? 46'b1100000010011110100111011000000100111101001110 :
(key == 11'b10111011101) ? 46'b1100000001111000010111011000000011110000101110 :
(key == 11'b10111011110) ? 46'b1100000001010010001010011000000010100100010100 :
(key == 11'b10111011111) ? 46'b1100000000101011111110111000000001010111111101 :
(key == 11'b10111100000) ? 46'b1100000000000101110110011000000000001011101100 :
(key == 11'b10111100001) ? 46'b1011111111011111101111010111111110111111011110 :
(key == 11'b10111100010) ? 46'b1011111110111001101011010111111101110011010110 :
(key == 11'b10111100011) ? 46'b1011111110010011101010010111111100100111010100 :
(key == 11'b10111100100) ? 46'b1011111101101101101011010111111011011011010110 :
(key == 11'b10111100101) ? 46'b1011111101000111101111010111111010001111011110 :
(key == 11'b10111100110) ? 46'b1011111100100001110100110111111001000011101001 :
(key == 11'b10111100111) ? 46'b1011111011111011111100110111110111110111111001 :
(key == 11'b10111101000) ? 46'b1011111011010110000111110111110110101100001111 :
(key == 11'b10111101001) ? 46'b1011111010110000010100010111110101100000101000 :
(key == 11'b10111101010) ? 46'b1011111010001010100011110111110100010101000111 :
(key == 11'b10111101011) ? 46'b1011111001100100110110010111110011001001101100 :
(key == 11'b10111101100) ? 46'b1011111000111111001010010111110001111110010100 :
(key == 11'b10111101101) ? 46'b1011111000011001100001010111110000110011000010 :
(key == 11'b10111101110) ? 46'b1011110111110011111001110111101111100111110011 :
(key == 11'b10111101111) ? 46'b1011110111001110010101010111101110011100101010 :
(key == 11'b10111110000) ? 46'b1011110110101000110010010111101101010001100100 :
(key == 11'b10111110001) ? 46'b1011110110000011010010010111101100000110100100 :
(key == 11'b10111110010) ? 46'b1011110101011101110101010111101010111011101010 :
(key == 11'b10111110011) ? 46'b1011110100111000011010010111101001110000110100 :
(key == 11'b10111110100) ? 46'b1011110100010011000001010111101000100110000010 :
(key == 11'b10111110101) ? 46'b1011110011101101101010010111100111011011010100 :
(key == 11'b10111110110) ? 46'b1011110011001000010110010111100110010000101100 :
(key == 11'b10111110111) ? 46'b1011110010100011000101010111100101000110001010 :
(key == 11'b10111111000) ? 46'b1011110001111101110101110111100011111011101011 :
(key == 11'b10111111001) ? 46'b1011110001011000101000010111100010110001010000 :
(key == 11'b10111111010) ? 46'b1011110000110011011101010111100001100110111010 :
(key == 11'b10111111011) ? 46'b1011110000001110010100110111100000011100101001 :
(key == 11'b10111111100) ? 46'b1011101111101001001111110111011111010010011111 :
(key == 11'b10111111101) ? 46'b1011101111000100001011010111011110001000010110 :
(key == 11'b10111111110) ? 46'b1011101110011111001010010111011100111110010100 :
(key == 11'b10111111111) ? 46'b1011101101111010001011010111011011110100010110 :
(key == 11'b11000000000) ? 46'b1011101101010101001101110111011010101010011011 :
(key == 11'b11000000001) ? 46'b1011101100110000010011010111011001100000100110 :
(key == 11'b11000000010) ? 46'b1011101100001011011011110111011000010110110111 :
(key == 11'b11000000011) ? 46'b1011101011100110100101110111010111001101001011 :
(key == 11'b11000000100) ? 46'b1011101011000001110001010111010110000011100010 :
(key == 11'b11000000101) ? 46'b1011101010011100111111110111010100111001111111 :
(key == 11'b11000000110) ? 46'b1011101001111000010001010111010011110000100010 :
(key == 11'b11000000111) ? 46'b1011101001010011100101010111010010100111001010 :
(key == 11'b11000001000) ? 46'b1011101000101110111010010111010001011101110100 :
(key == 11'b11000001001) ? 46'b1011101000001010010001110111010000010100100011 :
(key == 11'b11000001010) ? 46'b1011100111100101101100010111001111001011011000 :
(key == 11'b11000001011) ? 46'b1011100111000001001000010111001110000010010000 :
(key == 11'b11000001100) ? 46'b1011100110011100100111010111001100111001001110 :
(key == 11'b11000001101) ? 46'b1011100101111000000111110111001011110000001111 :
(key == 11'b11000001110) ? 46'b1011100101010011101011010111001010100111010110 :
(key == 11'b11000001111) ? 46'b1011100100101111010000010111001001011110100000 :
(key == 11'b11000010000) ? 46'b1011100100001010111000010111001000010101110000 :
(key == 11'b11000010001) ? 46'b1011100011100110100001110111000111001101000011 :
(key == 11'b11000010010) ? 46'b1011100011000010001110010111000110000100011100 :
(key == 11'b11000010011) ? 46'b1011100010011101111101010111000100111011111010 :
(key == 11'b11000010100) ? 46'b1011100001111001101101010111000011110011011010 :
(key == 11'b11000010101) ? 46'b1011100001010101011111110111000010101010111111 :
(key == 11'b11000010110) ? 46'b1011100000110001010101010111000001100010101010 :
(key == 11'b11000010111) ? 46'b1011100000001101001100010111000000011010011000 :
(key == 11'b11000011000) ? 46'b1011011111101001000110010110111111010010001100 :
(key == 11'b11000011001) ? 46'b1011011111000101000001110110111110001010000011 :
(key == 11'b11000011010) ? 46'b1011011110100000111111010110111101000001111110 :
(key == 11'b11000011011) ? 46'b1011011101111101000000010110111011111010000000 :
(key == 11'b11000011100) ? 46'b1011011101011001000010010110111010110010000100 :
(key == 11'b11000011101) ? 46'b1011011100110101000110010110111001101010001100 :
(key == 11'b11000011110) ? 46'b1011011100010001001101110110111000100010011011 :
(key == 11'b11000011111) ? 46'b1011011011101101010110110110110111011010101101 :
(key == 11'b11000100000) ? 46'b1011011011001001100010010110110110010011000100 :
(key == 11'b11000100001) ? 46'b1011011010100101101110110110110101001011011101 :
(key == 11'b11000100010) ? 46'b1011011010000001111110010110110100000011111100 :
(key == 11'b11000100011) ? 46'b1011011001011110001111110110110010111100011111 :
(key == 11'b11000100100) ? 46'b1011011000111010100100110110110001110101001001 :
(key == 11'b11000100101) ? 46'b1011011000010110111011010110110000101101110110 :
(key == 11'b11000100110) ? 46'b1011010111110011010011010110101111100110100110 :
(key == 11'b11000100111) ? 46'b1011010111001111101100110110101110011111011001 :
(key == 11'b11000101000) ? 46'b1011010110101100001010010110101101011000010100 :
(key == 11'b11000101001) ? 46'b1011010110001000101000110110101100010001010001 :
(key == 11'b11000101010) ? 46'b1011010101100101001001110110101011001010010011 :
(key == 11'b11000101011) ? 46'b1011010101000001101100010110101010000011011000 :
(key == 11'b11000101100) ? 46'b1011010100011110010001110110101000111100100011 :
(key == 11'b11000101101) ? 46'b1011010011111010111001010110100111110101110010 :
(key == 11'b11000101110) ? 46'b1011010011010111100010110110100110101111000101 :
(key == 11'b11000101111) ? 46'b1011010010110100001111010110100101101000011110 :
(key == 11'b11000110000) ? 46'b1011010010010000111100110110100100100001111001 :
(key == 11'b11000110001) ? 46'b1011010001101101101100110110100011011011011001 :
(key == 11'b11000110010) ? 46'b1011010001001010011111010110100010010100111110 :
(key == 11'b11000110011) ? 46'b1011010000100111010010110110100001001110100101 :
(key == 11'b11000110100) ? 46'b1011010000000100001001010110100000001000010010 :
(key == 11'b11000110101) ? 46'b1011001111100001000001110110011111000010000011 :
(key == 11'b11000110110) ? 46'b1011001110111101111100010110011101111011111000 :
(key == 11'b11000110111) ? 46'b1011001110011010111001010110011100110101110010 :
(key == 11'b11000111000) ? 46'b1011001101110111111000010110011011101111110000 :
(key == 11'b11000111001) ? 46'b1011001101010100111001010110011010101001110010 :
(key == 11'b11000111010) ? 46'b1011001100110001111100110110011001100011111001 :
(key == 11'b11000111011) ? 46'b1011001100001111000001110110011000011110000011 :
(key == 11'b11000111100) ? 46'b1011001011101100001000010110010111011000010000 :
(key == 11'b11000111101) ? 46'b1011001011001001010001110110010110010010100011 :
(key == 11'b11000111110) ? 46'b1011001010100110011101010110010101001100111010 :
(key == 11'b11000111111) ? 46'b1011001010000011101010110110010100000111010101 :
(key == 11'b11001000000) ? 46'b1011001001100000111010010110010011000001110100 :
(key == 11'b11001000001) ? 46'b1011001000111110001100110110010001111100011001 :
(key == 11'b11001000010) ? 46'b1011001000011011100000010110010000110111000000 :
(key == 11'b11001000011) ? 46'b1011000111111000110101010110001111110001101010 :
(key == 11'b11001000100) ? 46'b1011000111010110001101010110001110101100011010 :
(key == 11'b11001000101) ? 46'b1011000110110011100111010110001101100111001110 :
(key == 11'b11001000110) ? 46'b1011000110010001000100010110001100100010001000 :
(key == 11'b11001000111) ? 46'b1011000101101110100010010110001011011101000100 :
(key == 11'b11001001000) ? 46'b1011000101001100000010010110001010011000000100 :
(key == 11'b11001001001) ? 46'b1011000100101001100100010110001001010011001000 :
(key == 11'b11001001010) ? 46'b1011000100000111001000110110001000001110010001 :
(key == 11'b11001001011) ? 46'b1011000011100100101111010110000111001001011110 :
(key == 11'b11001001100) ? 46'b1011000011000010010111110110000110000100101111 :
(key == 11'b11001001101) ? 46'b1011000010100000000010010110000101000000000100 :
(key == 11'b11001001110) ? 46'b1011000001111101101111010110000011111011011110 :
(key == 11'b11001001111) ? 46'b1011000001011011011101010110000010110110111010 :
(key == 11'b11001010000) ? 46'b1011000000111001001101110110000001110010011011 :
(key == 11'b11001010001) ? 46'b1011000000010111000000010110000000101110000000 :
(key == 11'b11001010010) ? 46'b1010111111110100110100110101111111101001101001 :
(key == 11'b11001010011) ? 46'b1010111111010010101100010101111110100101011000 :
(key == 11'b11001010100) ? 46'b1010111110110000100100110101111101100001001001 :
(key == 11'b11001010101) ? 46'b1010111110001110011111110101111100011100111111 :
(key == 11'b11001010110) ? 46'b1010111101101100011100010101111011011000111000 :
(key == 11'b11001010111) ? 46'b1010111101001010011010010101111010010100110100 :
(key == 11'b11001011000) ? 46'b1010111100101000011011010101111001010000110110 :
(key == 11'b11001011001) ? 46'b1010111100000110011101110101111000001100111011 :
(key == 11'b11001011010) ? 46'b1010111011100100100011010101110111001001000110 :
(key == 11'b11001011011) ? 46'b1010111011000010101010010101110110000101010100 :
(key == 11'b11001011100) ? 46'b1010111010100000110010110101110101000001100101 :
(key == 11'b11001011101) ? 46'b1010111001111110111101010101110011111101111010 :
(key == 11'b11001011110) ? 46'b1010111001011101001001110101110010111010010011 :
(key == 11'b11001011111) ? 46'b1010111000111011011001010101110001110110110010 :
(key == 11'b11001100000) ? 46'b1010111000011001101001110101110000110011010011 :
(key == 11'b11001100001) ? 46'b1010110111110111111100110101101111101111111001 :
(key == 11'b11001100010) ? 46'b1010110111010110010001010101101110101100100010 :
(key == 11'b11001100011) ? 46'b1010110110110100100111010101101101101001001110 :
(key == 11'b11001100100) ? 46'b1010110110010011000000010101101100100110000000 :
(key == 11'b11001100101) ? 46'b1010110101110001011010110101101011100010110101 :
(key == 11'b11001100110) ? 46'b1010110101001111110111010101101010011111101110 :
(key == 11'b11001100111) ? 46'b1010110100101110010101110101101001011100101011 :
(key == 11'b11001101000) ? 46'b1010110100001100110110010101101000011001101100 :
(key == 11'b11001101001) ? 46'b1010110011101011011001010101100111010110110010 :
(key == 11'b11001101010) ? 46'b1010110011001001111101010101100110010011111010 :
(key == 11'b11001101011) ? 46'b1010110010101000100011110101100101010001000111 :
(key == 11'b11001101100) ? 46'b1010110010000111001100010101100100001110011000 :
(key == 11'b11001101101) ? 46'b1010110001100101110110110101100011001011101101 :
(key == 11'b11001101110) ? 46'b1010110001000100100011010101100010001001000110 :
(key == 11'b11001101111) ? 46'b1010110000100011010001010101100001000110100010 :
(key == 11'b11001110000) ? 46'b1010110000000010000000110101100000000100000001 :
(key == 11'b11001110001) ? 46'b1010101111100000110011010101011111000001100110 :
(key == 11'b11001110010) ? 46'b1010101110111111100111010101011101111111001110 :
(key == 11'b11001110011) ? 46'b1010101110011110011100110101011100111100111001 :
(key == 11'b11001110100) ? 46'b1010101101111101010101010101011011111010101010 :
(key == 11'b11001110101) ? 46'b1010101101011100001110010101011010111000011100 :
(key == 11'b11001110110) ? 46'b1010101100111011001010010101011001110110010100 :
(key == 11'b11001110111) ? 46'b1010101100011010000111110101011000110100001111 :
(key == 11'b11001111000) ? 46'b1010101011111001000111110101010111110010001111 :
(key == 11'b11001111001) ? 46'b1010101011011000001001010101010110110000010010 :
(key == 11'b11001111010) ? 46'b1010101010110111001100010101010101101110011000 :
(key == 11'b11001111011) ? 46'b1010101010010110010000110101010100101100100001 :
(key == 11'b11001111100) ? 46'b1010101001110101011000010101010011101010110000 :
(key == 11'b11001111101) ? 46'b1010101001010100100001010101010010101001000010 :
(key == 11'b11001111110) ? 46'b1010101000110011101100010101010001100111011000 :
(key == 11'b11001111111) ? 46'b1010101000010010111001010101010000100101110010 :
(key == 11'b11010000000) ? 46'b1010100111110010001000010101001111100100010000 :
(key == 11'b11010000001) ? 46'b1010100111010001011000110101001110100010110001 :
(key == 11'b11010000010) ? 46'b1010100110110000101010110101001101100001010101 :
(key == 11'b11010000011) ? 46'b1010100110001111111111010101001100011111111110 :
(key == 11'b11010000100) ? 46'b1010100101101111010100110101001011011110101001 :
(key == 11'b11010000101) ? 46'b1010100101001110101101010101001010011101011010 :
(key == 11'b11010000110) ? 46'b1010100100101110000111110101001001011100001111 :
(key == 11'b11010000111) ? 46'b1010100100001101100100010101001000011011001000 :
(key == 11'b11010001000) ? 46'b1010100011101101000001010101000111011010000010 :
(key == 11'b11010001001) ? 46'b1010100011001100100001010101000110011001000010 :
(key == 11'b11010001010) ? 46'b1010100010101100000010110101000101011000000101 :
(key == 11'b11010001011) ? 46'b1010100010001011100110010101000100010111001100 :
(key == 11'b11010001100) ? 46'b1010100001101011001010110101000011010110010101 :
(key == 11'b11010001101) ? 46'b1010100001001010110001110101000010010101100011 :
(key == 11'b11010001110) ? 46'b1010100000101010011011010101000001010100110110 :
(key == 11'b11010001111) ? 46'b1010100000001010000101110101000000010100001011 :
(key == 11'b11010010000) ? 46'b1010011111101001110010110100111111010011100101 :
(key == 11'b11010010001) ? 46'b1010011111001001100001010100111110010011000010 :
(key == 11'b11010010010) ? 46'b1010011110101001010001010100111101010010100010 :
(key == 11'b11010010011) ? 46'b1010011110001001000011010100111100010010000110 :
(key == 11'b11010010100) ? 46'b1010011101101000110111010100111011010001101110 :
(key == 11'b11010010101) ? 46'b1010011101001000101101010100111010010001011010 :
(key == 11'b11010010110) ? 46'b1010011100101000100100110100111001010001001001 :
(key == 11'b11010010111) ? 46'b1010011100001000011110010100111000010000111100 :
(key == 11'b11010011000) ? 46'b1010011011101000011001110100110111010000110011 :
(key == 11'b11010011001) ? 46'b1010011011001000010110010100110110010000101100 :
(key == 11'b11010011010) ? 46'b1010011010101000010101010100110101010000101010 :
(key == 11'b11010011011) ? 46'b1010011010001000010110110100110100010000101101 :
(key == 11'b11010011100) ? 46'b1010011001101000011000110100110011010000110001 :
(key == 11'b11010011101) ? 46'b1010011001001000011101110100110010010000111011 :
(key == 11'b11010011110) ? 46'b1010011000101000100011010100110001010001000110 :
(key == 11'b11010011111) ? 46'b1010011000001000101010110100110000010001010101 :
(key == 11'b11010100000) ? 46'b1010010111101000110101010100101111010001101010 :
(key == 11'b11010100001) ? 46'b1010010111001001000000110100101110010010000001 :
(key == 11'b11010100010) ? 46'b1010010110101001001110010100101101010010011100 :
(key == 11'b11010100011) ? 46'b1010010110001001011100110100101100010010111001 :
(key == 11'b11010100100) ? 46'b1010010101101001101101110100101011010011011011 :
(key == 11'b11010100101) ? 46'b1010010101001010000001010100101010010100000010 :
(key == 11'b11010100110) ? 46'b1010010100101010010101110100101001010100101011 :
(key == 11'b11010100111) ? 46'b1010010100001010101100010100101000010101011000 :
(key == 11'b11010101000) ? 46'b1010010011101011000011110100100111010110000111 :
(key == 11'b11010101001) ? 46'b1010010011001011011101110100100110010110111011 :
(key == 11'b11010101010) ? 46'b1010010010101011111010010100100101010111110100 :
(key == 11'b11010101011) ? 46'b1010010010001100010111110100100100011000101111 :
(key == 11'b11010101100) ? 46'b1010010001101100110110010100100011011001101100 :
(key == 11'b11010101101) ? 46'b1010010001001101010111110100100010011010101111 :
(key == 11'b11010101110) ? 46'b1010010000101101111010110100100001011011110101 :
(key == 11'b11010101111) ? 46'b1010010000001110011111010100100000011100111110 :
(key == 11'b11010110000) ? 46'b1010001111101111000101010100011111011110001010 :
(key == 11'b11010110001) ? 46'b1010001111001111101100110100011110011111011001 :
(key == 11'b11010110010) ? 46'b1010001110110000010111010100011101100000101110 :
(key == 11'b11010110011) ? 46'b1010001110010001000010010100011100100010000100 :
(key == 11'b11010110100) ? 46'b1010001101110001101111010100011011100011011110 :
(key == 11'b11010110101) ? 46'b1010001101010010011110010100011010100100111100 :
(key == 11'b11010110110) ? 46'b1010001100110011001111010100011001100110011110 :
(key == 11'b11010110111) ? 46'b1010001100010100000010010100011000101000000100 :
(key == 11'b11010111000) ? 46'b1010001011110100110110010100010111101001101100 :
(key == 11'b11010111001) ? 46'b1010001011010101101100010100010110101011011000 :
(key == 11'b11010111010) ? 46'b1010001010110110100100010100010101101101001000 :
(key == 11'b11010111011) ? 46'b1010001010010111011101110100010100101110111011 :
(key == 11'b11010111100) ? 46'b1010001001111000011000110100010011110000110001 :
(key == 11'b11010111101) ? 46'b1010001001011001010110010100010010110010101100 :
(key == 11'b11010111110) ? 46'b1010001000111010010100110100010001110100101001 :
(key == 11'b11010111111) ? 46'b1010001000011011010101110100010000110110101011 :
(key == 11'b11011000000) ? 46'b1010000111111100011000010100001111111000110000 :
(key == 11'b11011000001) ? 46'b1010000111011101011011010100001110111010110110 :
(key == 11'b11011000010) ? 46'b1010000110111110100000010100001101111101000000 :
(key == 11'b11011000011) ? 46'b1010000110011111101000010100001100111111010000 :
(key == 11'b11011000100) ? 46'b1010000110000000110001010100001100000001100010 :
(key == 11'b11011000101) ? 46'b1010000101100001111100010100001011000011111000 :
(key == 11'b11011000110) ? 46'b1010000101000011001000010100001010000110010000 :
(key == 11'b11011000111) ? 46'b1010000100100100010110110100001001001000101101 :
(key == 11'b11011001000) ? 46'b1010000100000101100110110100001000001011001101 :
(key == 11'b11011001001) ? 46'b1010000011100110111000010100000111001101110000 :
(key == 11'b11011001010) ? 46'b1010000011001000001011010100000110010000010110 :
(key == 11'b11011001011) ? 46'b1010000010101001011111110100000101010010111111 :
(key == 11'b11011001100) ? 46'b1010000010001010110110010100000100010101101100 :
(key == 11'b11011001101) ? 46'b1010000001101100001110110100000011011000011101 :
(key == 11'b11011001110) ? 46'b1010000001001101101001010100000010011011010010 :
(key == 11'b11011001111) ? 46'b1010000000101111000101010100000001011110001010 :
(key == 11'b11011010000) ? 46'b1010000000010000100010110100000000100001000101 :
(key == 11'b11011010001) ? 46'b1001111111110010000001110011111111100100000011 :
(key == 11'b11011010010) ? 46'b1001111111010011100010010011111110100111000100 :
(key == 11'b11011010011) ? 46'b1001111110110101000100010011111101101010001000 :
(key == 11'b11011010100) ? 46'b1001111110010110100111110011111100101101001111 :
(key == 11'b11011010101) ? 46'b1001111101111000001110010011111011110000011100 :
(key == 11'b11011010110) ? 46'b1001111101011001110101010011111010110011101010 :
(key == 11'b11011010111) ? 46'b1001111100111011011110010011111001110110111100 :
(key == 11'b11011011000) ? 46'b1001111100011101001001010011111000111010010010 :
(key == 11'b11011011001) ? 46'b1001111011111110110101110011110111111101101011 :
(key == 11'b11011011010) ? 46'b1001111011100000100011110011110111000001000111 :
(key == 11'b11011011011) ? 46'b1001111011000010010011010011110110000100100110 :
(key == 11'b11011011100) ? 46'b1001111010100100000100010011110101001000001000 :
(key == 11'b11011011101) ? 46'b1001111010000101110111010011110100001011101110 :
(key == 11'b11011011110) ? 46'b1001111001100111101100010011110011001111011000 :
(key == 11'b11011011111) ? 46'b1001111001001001100011010011110010010011000110 :
(key == 11'b11011100000) ? 46'b1001111000101011011011010011110001010110110110 :
(key == 11'b11011100001) ? 46'b1001111000001101010100010011110000011010101000 :
(key == 11'b11011100010) ? 46'b1001110111101111001111110011101111011110011111 :
(key == 11'b11011100011) ? 46'b1001110111010001001100110011101110100010011001 :
(key == 11'b11011100100) ? 46'b1001110110110011001011010011101101100110010110 :
(key == 11'b11011100101) ? 46'b1001110110010101001011010011101100101010010110 :
(key == 11'b11011100110) ? 46'b1001110101110111001100110011101011101110011001 :
(key == 11'b11011100111) ? 46'b1001110101011001001111110011101010110010011111 :
(key == 11'b11011101000) ? 46'b1001110100111011010101010011101001110110101010 :
(key == 11'b11011101001) ? 46'b1001110100011101011011110011101000111010110111 :
(key == 11'b11011101010) ? 46'b1001110011111111100100010011100111111111001000 :
(key == 11'b11011101011) ? 46'b1001110011100001101101110011100111000011011011 :
(key == 11'b11011101100) ? 46'b1001110011000011111001110011100110000111110011 :
(key == 11'b11011101101) ? 46'b1001110010100110000111010011100101001100001110 :
(key == 11'b11011101110) ? 46'b1001110010001000010101010011100100010000101010 :
(key == 11'b11011101111) ? 46'b1001110001101010100101010011100011010101001010 :
(key == 11'b11011110000) ? 46'b1001110001001100110111010011100010011001101110 :
(key == 11'b11011110001) ? 46'b1001110000101111001010110011100001011110010101 :
(key == 11'b11011110010) ? 46'b1001110000010001100000010011100000100011000000 :
(key == 11'b11011110011) ? 46'b1001101111110011110111110011011111100111101111 :
(key == 11'b11011110100) ? 46'b1001101111010110001111110011011110101100011111 :
(key == 11'b11011110101) ? 46'b1001101110111000101001010011011101110001010010 :
(key == 11'b11011110110) ? 46'b1001101110011011000101010011011100110110001010 :
(key == 11'b11011110111) ? 46'b1001101101111101100010010011011011111011000100 :
(key == 11'b11011111000) ? 46'b1001101101100000000001010011011011000000000010 :
(key == 11'b11011111001) ? 46'b1001101101000010100001010011011010000101000010 :
(key == 11'b11011111010) ? 46'b1001101100100101000011010011011001001010000110 :
(key == 11'b11011111011) ? 46'b1001101100000111100110010011011000001111001100 :
(key == 11'b11011111100) ? 46'b1001101011101010001011110011010111010100010111 :
(key == 11'b11011111101) ? 46'b1001101011001100110010110011010110011001100101 :
(key == 11'b11011111110) ? 46'b1001101010101111011010010011010101011110110100 :
(key == 11'b11011111111) ? 46'b1001101010010010000011110011010100100100000111 :
(key == 11'b11100000000) ? 46'b1001101001110100101111010011010011101001011110 :
(key == 11'b11100000001) ? 46'b1001101001010111011100010011010010101110111000 :
(key == 11'b11100000010) ? 46'b1001101000111010001010110011010001110100010101 :
(key == 11'b11100000011) ? 46'b1001101000011100111010110011010000111001110101 :
(key == 11'b11100000100) ? 46'b1001100111111111101101010011001111111111011010 :
(key == 11'b11100000101) ? 46'b1001100111100010100000110011001111000101000001 :
(key == 11'b11100000110) ? 46'b1001100111000101010101010011001110001010101010 :
(key == 11'b11100000111) ? 46'b1001100110101000001011010011001101010000010110 :
(key == 11'b11100001000) ? 46'b1001100110001011000010110011001100010110000101 :
(key == 11'b11100001001) ? 46'b1001100101101101111011110011001011011011110111 :
(key == 11'b11100001010) ? 46'b1001100101010000110111010011001010100001101110 :
(key == 11'b11100001011) ? 46'b1001100100110011110011110011001001100111100111 :
(key == 11'b11100001100) ? 46'b1001100100010110110010010011001000101101100100 :
(key == 11'b11100001101) ? 46'b1001100011111001110001110011000111110011100011 :
(key == 11'b11100001110) ? 46'b1001100011011100110010010011000110111001100100 :
(key == 11'b11100001111) ? 46'b1001100010111111110101010011000101111111101010 :
(key == 11'b11100010000) ? 46'b1001100010100010111001010011000101000101110010 :
(key == 11'b11100010001) ? 46'b1001100010000101111111110011000100001011111111 :
(key == 11'b11100010010) ? 46'b1001100001101001000110010011000011010010001100 :
(key == 11'b11100010011) ? 46'b1001100001001100001111110011000010011000011111 :
(key == 11'b11100010100) ? 46'b1001100000101111011010010011000001011110110100 :
(key == 11'b11100010101) ? 46'b1001100000010010100101110011000000100101001011 :
(key == 11'b11100010110) ? 46'b1001011111110101110011010010111111101011100110 :
(key == 11'b11100010111) ? 46'b1001011111011001000001110010111110110010000011 :
(key == 11'b11100011000) ? 46'b1001011110111100010010110010111101111000100101 :
(key == 11'b11100011001) ? 46'b1001011110011111100100010010111100111111001000 :
(key == 11'b11100011010) ? 46'b1001011110000010110111110010111100000101101111 :
(key == 11'b11100011011) ? 46'b1001011101100110001101010010111011001100011010 :
(key == 11'b11100011100) ? 46'b1001011101001001100011010010111010010011000110 :
(key == 11'b11100011101) ? 46'b1001011100101100111011010010111001011001110110 :
(key == 11'b11100011110) ? 46'b1001011100010000010101010010111000100000101010 :
(key == 11'b11100011111) ? 46'b1001011011110011110000010010110111100111100000 :
(key == 11'b11100100000) ? 46'b1001011011010111001100010010110110101110011000 :
(key == 11'b11100100001) ? 46'b1001011010111010101010110010110101110101010101 :
(key == 11'b11100100010) ? 46'b1001011010011110001010010010110100111100010100 :
(key == 11'b11100100011) ? 46'b1001011010000001101010110010110100000011010101 :
(key == 11'b11100100100) ? 46'b1001011001100101001101110010110011001010011011 :
(key == 11'b11100100101) ? 46'b1001011001001000110010010010110010010001100100 :
(key == 11'b11100100110) ? 46'b1001011000101100010111010010110001011000101110 :
(key == 11'b11100100111) ? 46'b1001011000001111111110010010110000011111111100 :
(key == 11'b11100101000) ? 46'b1001010111110011100111010010101111100111001110 :
(key == 11'b11100101001) ? 46'b1001010111010111010001010010101110101110100010 :
(key == 11'b11100101010) ? 46'b1001010110111010111100010010101101110101111000 :
(key == 11'b11100101011) ? 46'b1001010110011110101001010010101100111101010010 :
(key == 11'b11100101100) ? 46'b1001010110000010010111010010101100000100101110 :
(key == 11'b11100101101) ? 46'b1001010101100110000111110010101011001100001111 :
(key == 11'b11100101110) ? 46'b1001010101001001111001010010101010010011110010 :
(key == 11'b11100101111) ? 46'b1001010100101101101011110010101001011011010111 :
(key == 11'b11100110000) ? 46'b1001010100010001100000010010101000100011000000 :
(key == 11'b11100110001) ? 46'b1001010011110101010101110010100111101010101011 :
(key == 11'b11100110010) ? 46'b1001010011011001001101010010100110110010011010 :
(key == 11'b11100110011) ? 46'b1001010010111101000101110010100101111010001011 :
(key == 11'b11100110100) ? 46'b1001010010100001000000010010100101000010000000 :
(key == 11'b11100110101) ? 46'b1001010010000100111011110010100100001001110111 :
(key == 11'b11100110110) ? 46'b1001010001101000111000010010100011010001110000 :
(key == 11'b11100110111) ? 46'b1001010001001100110111010010100010011001101110 :
(key == 11'b11100111000) ? 46'b1001010000110000110111010010100001100001101110 :
(key == 11'b11100111001) ? 46'b1001010000010100111000010010100000101001110000 :
(key == 11'b11100111010) ? 46'b1001001111111000111011010010011111110001110110 :
(key == 11'b11100111011) ? 46'b1001001111011101000000010010011110111010000000 :
(key == 11'b11100111100) ? 46'b1001001111000001000101110010011110000010001011 :
(key == 11'b11100111101) ? 46'b1001001110100101001100110010011101001010011001 :
(key == 11'b11100111110) ? 46'b1001001110001001010101010010011100010010101010 :
(key == 11'b11100111111) ? 46'b1001001101101101011111010010011011011010111110 :
(key == 11'b11101000000) ? 46'b1001001101010001101011010010011010100011010110 :
(key == 11'b11101000001) ? 46'b1001001100110101111001010010011001101011110010 :
(key == 11'b11101000010) ? 46'b1001001100011010000111010010011000110100001110 :
(key == 11'b11101000011) ? 46'b1001001011111110010110010010010111111100101100 :
(key == 11'b11101000100) ? 46'b1001001011100010100111110010010111000101001111 :
(key == 11'b11101000101) ? 46'b1001001011000110111010110010010110001101110101 :
(key == 11'b11101000110) ? 46'b1001001010101011001111010010010101010110011110 :
(key == 11'b11101000111) ? 46'b1001001010001111100101010010010100011111001010 :
(key == 11'b11101001000) ? 46'b1001001001110011111100010010010011100111111000 :
(key == 11'b11101001001) ? 46'b1001001001011000010100010010010010110000101000 :
(key == 11'b11101001010) ? 46'b1001001000111100101110110010010001111001011101 :
(key == 11'b11101001011) ? 46'b1001001000100001001001010010010001000010010010 :
(key == 11'b11101001100) ? 46'b1001001000000101100110110010010000001011001101 :
(key == 11'b11101001101) ? 46'b1001000111101010000100010010001111010100001000 :
(key == 11'b11101001110) ? 46'b1001000111001110100100010010001110011101001000 :
(key == 11'b11101001111) ? 46'b1001000110110011000101010010001101100110001010 :
(key == 11'b11101010000) ? 46'b1001000110010111100111010010001100101111001110 :
(key == 11'b11101010001) ? 46'b1001000101111100001010110010001011111000010101 :
(key == 11'b11101010010) ? 46'b1001000101100000101111110010001011000001011111 :
(key == 11'b11101010011) ? 46'b1001000101000101010110010010001010001010101100 :
(key == 11'b11101010100) ? 46'b1001000100101001111110010010001001010011111100 :
(key == 11'b11101010101) ? 46'b1001000100001110100111110010001000011101001111 :
(key == 11'b11101010110) ? 46'b1001000011110011010010110010000111100110100101 :
(key == 11'b11101010111) ? 46'b1001000011010111111111010010000110101111111110 :
(key == 11'b11101011000) ? 46'b1001000010111100101101010010000101111001011010 :
(key == 11'b11101011001) ? 46'b1001000010100001011100010010000101000010111000 :
(key == 11'b11101011010) ? 46'b1001000010000110001100010010000100001100011000 :
(key == 11'b11101011011) ? 46'b1001000001101010111110010010000011010101111100 :
(key == 11'b11101011100) ? 46'b1001000001001111110001010010000010011111100010 :
(key == 11'b11101011101) ? 46'b1001000000110100100101010010000001101001001010 :
(key == 11'b11101011110) ? 46'b1001000000011001011010110010000000110010110101 :
(key == 11'b11101011111) ? 46'b1000111111111110010010010001111111111100100100 :
(key == 11'b11101100000) ? 46'b1000111111100011001011110001111111000110010111 :
(key == 11'b11101100001) ? 46'b1000111111001000000101110001111110010000001011 :
(key == 11'b11101100010) ? 46'b1000111110101101000001010001111101011010000010 :
(key == 11'b11101100011) ? 46'b1000111110010001111110010001111100100011111100 :
(key == 11'b11101100100) ? 46'b1000111101110110111100010001111011101101111000 :
(key == 11'b11101100101) ? 46'b1000111101011011111011010001111010110111110110 :
(key == 11'b11101100110) ? 46'b1000111101000000111100010001111010000001111000 :
(key == 11'b11101100111) ? 46'b1000111100100101111110010001111001001011111100 :
(key == 11'b11101101000) ? 46'b1000111100001011000010010001111000010110000100 :
(key == 11'b11101101001) ? 46'b1000111011110000000111010001110111100000001110 :
(key == 11'b11101101010) ? 46'b1000111011010101001101010001110110101010011010 :
(key == 11'b11101101011) ? 46'b1000111010111010010100110001110101110100101001 :
(key == 11'b11101101100) ? 46'b1000111010011111011101110001110100111110111011 :
(key == 11'b11101101101) ? 46'b1000111010000100101000010001110100001001010000 :
(key == 11'b11101101110) ? 46'b1000111001101001110100010001110011010011101000 :
(key == 11'b11101101111) ? 46'b1000111001001111000001110001110010011110000011 :
(key == 11'b11101110000) ? 46'b1000111000110100010000010001110001101000100000 :
(key == 11'b11101110001) ? 46'b1000111000011001011111110001110000110010111111 :
(key == 11'b11101110010) ? 46'b1000110111111110110001010001101111111101100010 :
(key == 11'b11101110011) ? 46'b1000110111100100000011110001101111001000000111 :
(key == 11'b11101110100) ? 46'b1000110111001001010111010001101110010010101110 :
(key == 11'b11101110101) ? 46'b1000110110101110101100010001101101011101011000 :
(key == 11'b11101110110) ? 46'b1000110110010100000010110001101100101000000101 :
(key == 11'b11101110111) ? 46'b1000110101111001011010110001101011110010110101 :
(key == 11'b11101111000) ? 46'b1000110101011110110100010001101010111101101000 :
(key == 11'b11101111001) ? 46'b1000110101000100001111010001101010001000011110 :
(key == 11'b11101111010) ? 46'b1000110100101001101011010001101001010011010110 :
(key == 11'b11101111011) ? 46'b1000110100001111001000010001101000011110010000 :
(key == 11'b11101111100) ? 46'b1000110011110100100110010001100111101001001100 :
(key == 11'b11101111101) ? 46'b1000110011011010000110010001100110110100001100 :
(key == 11'b11101111110) ? 46'b1000110010111111101000010001100101111111010000 :
(key == 11'b11101111111) ? 46'b1000110010100101001010110001100101001010010101 :
(key == 11'b11110000000) ? 46'b1000110010001010101110110001100100010101011101 :
(key == 11'b11110000001) ? 46'b1000110001110000010011010001100011100000100110 :
(key == 11'b11110000010) ? 46'b1000110001010101111001110001100010101011110011 :
(key == 11'b11110000011) ? 46'b1000110000111011100001010001100001110111000010 :
(key == 11'b11110000100) ? 46'b1000110000100001001010110001100001000010010101 :
(key == 11'b11110000101) ? 46'b1000110000000110110101010001100000001101101010 :
(key == 11'b11110000110) ? 46'b1000101111101100100001110001011111011001000011 :
(key == 11'b11110000111) ? 46'b1000101111010010001110110001011110100100011101 :
(key == 11'b11110001000) ? 46'b1000101110110111111101010001011101101111111010 :
(key == 11'b11110001001) ? 46'b1000101110011101101100010001011100111011011000 :
(key == 11'b11110001010) ? 46'b1000101110000011011101010001011100000110111010 :
(key == 11'b11110001011) ? 46'b1000101101101001001111010001011011010010011110 :
(key == 11'b11110001100) ? 46'b1000101101001111000011010001011010011110000110 :
(key == 11'b11110001101) ? 46'b1000101100110100110111110001011001101001101111 :
(key == 11'b11110001110) ? 46'b1000101100011010101101110001011000110101011011 :
(key == 11'b11110001111) ? 46'b1000101100000000100110010001011000000001001100 :
(key == 11'b11110010000) ? 46'b1000101011100110011111010001010111001100111110 :
(key == 11'b11110010001) ? 46'b1000101011001100011000110001010110011000110001 :
(key == 11'b11110010010) ? 46'b1000101010110010010100010001010101100100101000 :
(key == 11'b11110010011) ? 46'b1000101010011000010000110001010100110000100001 :
(key == 11'b11110010100) ? 46'b1000101001111110001110010001010011111100011100 :
(key == 11'b11110010101) ? 46'b1000101001100100001110010001010011001000011100 :
(key == 11'b11110010110) ? 46'b1000101001001010001111010001010010010100011110 :
(key == 11'b11110010111) ? 46'b1000101000110000010000010001010001100000100000 :
(key == 11'b11110011000) ? 46'b1000101000010110010011010001010000101100100110 :
(key == 11'b11110011001) ? 46'b1000100111111100011000010001001111111000110000 :
(key == 11'b11110011010) ? 46'b1000100111100010011101010001001111000100111010 :
(key == 11'b11110011011) ? 46'b1000100111001000100100010001001110010001001000 :
(key == 11'b11110011100) ? 46'b1000100110101110101101010001001101011101011010 :
(key == 11'b11110011101) ? 46'b1000100110010100110110110001001100101001101101 :
(key == 11'b11110011110) ? 46'b1000100101111011000001010001001011110110000010 :
(key == 11'b11110011111) ? 46'b1000100101100001001100110001001011000010011001 :
(key == 11'b11110100000) ? 46'b1000100101000111011010010001001010001110110100 :
(key == 11'b11110100001) ? 46'b1000100100101101101000110001001001011011010001 :
(key == 11'b11110100010) ? 46'b1000100100010011111001010001001000100111110010 :
(key == 11'b11110100011) ? 46'b1000100011111010001010010001000111110100010100 :
(key == 11'b11110100100) ? 46'b1000100011100000011011110001000111000000110111 :
(key == 11'b11110100101) ? 46'b1000100011000110101111110001000110001101011111 :
(key == 11'b11110100110) ? 46'b1000100010101101000101010001000101011010001010 :
(key == 11'b11110100111) ? 46'b1000100010010011011010110001000100100110110101 :
(key == 11'b11110101000) ? 46'b1000100001111001110001110001000011110011100011 :
(key == 11'b11110101001) ? 46'b1000100001100000001011010001000011000000010110 :
(key == 11'b11110101010) ? 46'b1000100001000110100101010001000010001101001010 :
(key == 11'b11110101011) ? 46'b1000100000101100111111110001000001011001111111 :
(key == 11'b11110101100) ? 46'b1000100000010011011100110001000000100110111001 :
(key == 11'b11110101101) ? 46'b1000011111111001111001110000111111110011110011 :
(key == 11'b11110101110) ? 46'b1000011111100000011001010000111111000000110010 :
(key == 11'b11110101111) ? 46'b1000011111000110111001110000111110001101110011 :
(key == 11'b11110110000) ? 46'b1000011110101101011010010000111101011010110100 :
(key == 11'b11110110001) ? 46'b1000011110010011111100110000111100100111111001 :
(key == 11'b11110110010) ? 46'b1000011101111010100001010000111011110101000010 :
(key == 11'b11110110011) ? 46'b1000011101100001000110010000111011000010001100 :
(key == 11'b11110110100) ? 46'b1000011101000111101101010000111010001111011010 :
(key == 11'b11110110101) ? 46'b1000011100101110010100110000111001011100101001 :
(key == 11'b11110110110) ? 46'b1000011100010100111101010000111000101001111010 :
(key == 11'b11110110111) ? 46'b1000011011111011100110110000110111110111001101 :
(key == 11'b11110111000) ? 46'b1000011011100010010010110000110111000100100101 :
(key == 11'b11110111001) ? 46'b1000011011001000111110110000110110010001111101 :
(key == 11'b11110111010) ? 46'b1000011010101111101100010000110101011111011000 :
(key == 11'b11110111011) ? 46'b1000011010010110011011010000110100101100110110 :
(key == 11'b11110111100) ? 46'b1000011001111101001011110000110011111010010111 :
(key == 11'b11110111101) ? 46'b1000011001100011111101010000110011000111111010 :
(key == 11'b11110111110) ? 46'b1000011001001010101111110000110010010101011111 :
(key == 11'b11110111111) ? 46'b1000011000110001100011010000110001100011000110 :
(key == 11'b11111000000) ? 46'b1000011000011000011000010000110000110000110000 :
(key == 11'b11111000001) ? 46'b1000010111111111001110110000101111111110011101 :
(key == 11'b11111000010) ? 46'b1000010111100110000110110000101111001100001101 :
(key == 11'b11111000011) ? 46'b1000010111001100111111010000101110011001111110 :
(key == 11'b11111000100) ? 46'b1000010110110011111001110000101101100111110011 :
(key == 11'b11111000101) ? 46'b1000010110011010110100110000101100110101101001 :
(key == 11'b11111000110) ? 46'b1000010110000001110001010000101100000011100010 :
(key == 11'b11111000111) ? 46'b1000010101101000101110010000101011010001011100 :
(key == 11'b11111001000) ? 46'b1000010101001111101101010000101010011111011010 :
(key == 11'b11111001001) ? 46'b1000010100110110101100110000101001101101011001 :
(key == 11'b11111001010) ? 46'b1000010100011101101101110000101000111011011011 :
(key == 11'b11111001011) ? 46'b1000010100000100110000010000101000001001100000 :
(key == 11'b11111001100) ? 46'b1000010011101011110100010000100111010111101000 :
(key == 11'b11111001101) ? 46'b1000010011010010111001010000100110100101110010 :
(key == 11'b11111001110) ? 46'b1000010010111001111111010000100101110011111110 :
(key == 11'b11111001111) ? 46'b1000010010100001000110010000100101000010001100 :
(key == 11'b11111010000) ? 46'b1000010010001000001110110000100100010000011101 :
(key == 11'b11111010001) ? 46'b1000010001101111011000010000100011011110110000 :
(key == 11'b11111010010) ? 46'b1000010001010110100010110000100010101101000101 :
(key == 11'b11111010011) ? 46'b1000010000111101101111010000100001111011011110 :
(key == 11'b11111010100) ? 46'b1000010000100100111100010000100001001001111000 :
(key == 11'b11111010101) ? 46'b1000010000001100001001110000100000011000010011 :
(key == 11'b11111010110) ? 46'b1000001111110011011001110000011111100110110011 :
(key == 11'b11111010111) ? 46'b1000001111011010101010010000011110110101010100 :
(key == 11'b11111011000) ? 46'b1000001111000001111100110000011110000011111001 :
(key == 11'b11111011001) ? 46'b1000001110101001001111110000011101010010011111 :
(key == 11'b11111011010) ? 46'b1000001110010000100100010000011100100001001000 :
(key == 11'b11111011011) ? 46'b1000001101110111111001010000011011101111110010 :
(key == 11'b11111011100) ? 46'b1000001101011111010000010000011010111110100000 :
(key == 11'b11111011101) ? 46'b1000001101000110100111110000011010001101001111 :
(key == 11'b11111011110) ? 46'b1000001100101110000000110000011001011100000001 :
(key == 11'b11111011111) ? 46'b1000001100010101011010010000011000101010110100 :
(key == 11'b11111100000) ? 46'b1000001011111100110101110000010111111001101011 :
(key == 11'b11111100001) ? 46'b1000001011100100010001110000010111001000100011 :
(key == 11'b11111100010) ? 46'b1000001011001011110000010000010110010111100000 :
(key == 11'b11111100011) ? 46'b1000001010110011001111010000010101100110011110 :
(key == 11'b11111100100) ? 46'b1000001010011010101110110000010100110101011101 :
(key == 11'b11111100101) ? 46'b1000001010000010001111010000010100000100011110 :
(key == 11'b11111100110) ? 46'b1000001001101001110001010000010011010011100010 :
(key == 11'b11111100111) ? 46'b1000001001010001010100110000010010100010101001 :
(key == 11'b11111101000) ? 46'b1000001000111000111001110000010001110001110011 :
(key == 11'b11111101001) ? 46'b1000001000100000100000010000010001000001000000 :
(key == 11'b11111101010) ? 46'b1000001000001000000110110000010000010000001101 :
(key == 11'b11111101011) ? 46'b1000000111101111101110110000001111011111011101 :
(key == 11'b11111101100) ? 46'b1000000111010111011000010000001110101110110000 :
(key == 11'b11111101101) ? 46'b1000000110111111000010010000001101111110000100 :
(key == 11'b11111101110) ? 46'b1000000110100110101110010000001101001101011100 :
(key == 11'b11111101111) ? 46'b1000000110001110011010110000001100011100110101 :
(key == 11'b11111110000) ? 46'b1000000101110110001000110000001011101100010001 :
(key == 11'b11111110001) ? 46'b1000000101011101110111010000001010111011101110 :
(key == 11'b11111110010) ? 46'b1000000101000101100111110000001010001011001111 :
(key == 11'b11111110011) ? 46'b1000000100101101011000110000001001011010110001 :
(key == 11'b11111110100) ? 46'b1000000100010101001011010000001000101010010110 :
(key == 11'b11111110101) ? 46'b1000000011111100111110010000000111111001111100 :
(key == 11'b11111110110) ? 46'b1000000011100100110011010000000111001001100110 :
(key == 11'b11111110111) ? 46'b1000000011001100101000110000000110011001010001 :
(key == 11'b11111111000) ? 46'b1000000010110100011111110000000101101000111111 :
(key == 11'b11111111001) ? 46'b1000000010011100011000010000000100111000110000 :
(key == 11'b11111111010) ? 46'b1000000010000100010001010000000100001000100010 :
(key == 11'b11111111011) ? 46'b1000000001101100001100010000000011011000011000 :
(key == 11'b11111111100) ? 46'b1000000001010100000111110000000010101000001111 :
(key == 11'b11111111101) ? 46'b1000000000111100000100010000000001111000001000 :
(key == 11'b11111111110) ? 46'b1000000000100100000001110000000001001000000011 :
(key == 11'b11111111111) ? 46'b1000000000001100000000010000000000011000000000 : 46'd0;

endmodule

`default_nettype wire
