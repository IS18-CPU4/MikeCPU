`default_nettype none

module fsqrt_inv
   ( input wire [31:0] x,
     output wire [31:0] y,
     output wire ovf);

   // split sequence to each subsequence
   wire xs;
   wire [7:0] xe;
   wire [22:0] xm;
   assign {xs, xe, xm} = x;

   // calc s
   wire s;
   assign s = xs;

   wire [7:0] shift_xe;
   assign shift_xe = xe >> 1;

   // calc e
   wire [7:0] e;
   assign e = (xe[0] == 1) ? 8'd189 - shift_xe : 8'd190 - shift_xe; 

   // calc m
   wire [22:0] m;
   wire [47:0] val;
   wire [10:0] key;
   assign key = {xe[0], xm[22:13]};

   // lookup table and get constant and grad
   lookup_table lt(key, val);

   wire [24:0] constant;
   wire [22:0] grad;
   assign constant = val[47:23];
   assign grad = val[22:0];

   wire [47:0] grad2;
   assign grad2 = {1'b1, xm} * {1'b1, grad};

   wire [24:0] grad3;
   assign grad3 = (grad2[47] == 1'b0) ? {2'd0, grad2[46:24]} : {2'd0, grad2[47:25]};

   wire [24:0] tmp_m;
   assign tmp_m = constant - grad3;

   assign m = tmp_m[22:0]; // ignore implicit 1

   assign y = {s, e, m};
   assign ovf = 0;

endmodule

module lookup_table
   ( input wire [10:0] key,
     output wire [47:0] value);

   assign value =
(key == 11'b00000000000) ? 48'b100001111011101100111100000001111011101100111100 :
(key == 11'b00000000001) ? 48'b100001111010101001001010000001111010101001001010 :
(key == 11'b00000000010) ? 48'b100001111001100101011110000001111001100101011110 :
(key == 11'b00000000011) ? 48'b100001111000100001111000000001111000100001111000 :
(key == 11'b00000000100) ? 48'b100001110111011110011010000001110111011110011010 :
(key == 11'b00000000101) ? 48'b100001110110011011000001000001110110011011000001 :
(key == 11'b00000000110) ? 48'b100001110101010111101110000001110101010111101110 :
(key == 11'b00000000111) ? 48'b100001110100010100100010000001110100010100100010 :
(key == 11'b00000001000) ? 48'b100001110011010001011100000001110011010001011100 :
(key == 11'b00000001001) ? 48'b100001110010001110011100000001110010001110011100 :
(key == 11'b00000001010) ? 48'b100001110001001011100010000001110001001011100010 :
(key == 11'b00000001011) ? 48'b100001110000001000101111000001110000001000101111 :
(key == 11'b00000001100) ? 48'b100001101111000110000010000001101111000110000010 :
(key == 11'b00000001101) ? 48'b100001101110000011011100000001101110000011011100 :
(key == 11'b00000001110) ? 48'b100001101101000000111010000001101101000000111010 :
(key == 11'b00000001111) ? 48'b100001101011111110011111000001101011111110011111 :
(key == 11'b00000010000) ? 48'b100001101010111100001010000001101010111100001010 :
(key == 11'b00000010001) ? 48'b100001101001111001111100000001101001111001111100 :
(key == 11'b00000010010) ? 48'b100001101000110111110100000001101000110111110100 :
(key == 11'b00000010011) ? 48'b100001100111110101110010000001100111110101110010 :
(key == 11'b00000010100) ? 48'b100001100110110011110110000001100110110011110110 :
(key == 11'b00000010101) ? 48'b100001100101110001111111000001100101110001111111 :
(key == 11'b00000010110) ? 48'b100001100100110000001110000001100100110000001110 :
(key == 11'b00000010111) ? 48'b100001100011101110100100000001100011101110100100 :
(key == 11'b00000011000) ? 48'b100001100010101101000000000001100010101101000000 :
(key == 11'b00000011001) ? 48'b100001100001101011100011000001100001101011100011 :
(key == 11'b00000011010) ? 48'b100001100000101010001011000001100000101010001011 :
(key == 11'b00000011011) ? 48'b100001011111101000111000000001011111101000111000 :
(key == 11'b00000011100) ? 48'b100001011110100111101100000001011110100111101100 :
(key == 11'b00000011101) ? 48'b100001011101100110100101000001011101100110100101 :
(key == 11'b00000011110) ? 48'b100001011100100101100110000001011100100101100110 :
(key == 11'b00000011111) ? 48'b100001011011100100101011000001011011100100101011 :
(key == 11'b00000100000) ? 48'b100001011010100011110110000001011010100011110110 :
(key == 11'b00000100001) ? 48'b100001011001100011001000000001011001100011001000 :
(key == 11'b00000100010) ? 48'b100001011000100010011111000001011000100010011111 :
(key == 11'b00000100011) ? 48'b100001010111100001111101000001010111100001111101 :
(key == 11'b00000100100) ? 48'b100001010110100001100000000001010110100001100000 :
(key == 11'b00000100101) ? 48'b100001010101100001001000000001010101100001001000 :
(key == 11'b00000100110) ? 48'b100001010100100000110111000001010100100000110111 :
(key == 11'b00000100111) ? 48'b100001010011100000101100000001010011100000101100 :
(key == 11'b00000101000) ? 48'b100001010010100000100101000001010010100000100101 :
(key == 11'b00000101001) ? 48'b100001010001100000100101000001010001100000100101 :
(key == 11'b00000101010) ? 48'b100001010000100000101011000001010000100000101011 :
(key == 11'b00000101011) ? 48'b100001001111100000110110000001001111100000110110 :
(key == 11'b00000101100) ? 48'b100001001110100001001000000001001110100001001000 :
(key == 11'b00000101101) ? 48'b100001001101100001011110000001001101100001011110 :
(key == 11'b00000101110) ? 48'b100001001100100001111100000001001100100001111100 :
(key == 11'b00000101111) ? 48'b100001001011100010011110000001001011100010011110 :
(key == 11'b00000110000) ? 48'b100001001010100011000110000001001010100011000110 :
(key == 11'b00000110001) ? 48'b100001001001100011110011000001001001100011110011 :
(key == 11'b00000110010) ? 48'b100001001000100100100111000001001000100100100111 :
(key == 11'b00000110011) ? 48'b100001000111100101100000000001000111100101100000 :
(key == 11'b00000110100) ? 48'b100001000110100110011110000001000110100110011110 :
(key == 11'b00000110101) ? 48'b100001000101100111100011000001000101100111100011 :
(key == 11'b00000110110) ? 48'b100001000100101000101101000001000100101000101101 :
(key == 11'b00000110111) ? 48'b100001000011101001111100000001000011101001111100 :
(key == 11'b00000111000) ? 48'b100001000010101011010000000001000010101011010000 :
(key == 11'b00000111001) ? 48'b100001000001101100101100000001000001101100101100 :
(key == 11'b00000111010) ? 48'b100001000000101110001100000001000000101110001100 :
(key == 11'b00000111011) ? 48'b100000111111101111110001000000111111101111110001 :
(key == 11'b00000111100) ? 48'b100000111110110001011101000000111110110001011101 :
(key == 11'b00000111101) ? 48'b100000111101110011001110000000111101110011001110 :
(key == 11'b00000111110) ? 48'b100000111100110101000100000000111100110101000100 :
(key == 11'b00000111111) ? 48'b100000111011110111000000000000111011110111000000 :
(key == 11'b00001000000) ? 48'b100000111010111001000001000000111010111001000001 :
(key == 11'b00001000001) ? 48'b100000111001111011000111000000111001111011000111 :
(key == 11'b00001000010) ? 48'b100000111000111101010011000000111000111101010011 :
(key == 11'b00001000011) ? 48'b100000110111111111100110000000110111111111100110 :
(key == 11'b00001000100) ? 48'b100000110111000001111100000000110111000001111100 :
(key == 11'b00001000101) ? 48'b100000110110000100011000000000110110000100011000 :
(key == 11'b00001000110) ? 48'b100000110101000110111010000000110101000110111010 :
(key == 11'b00001000111) ? 48'b100000110100001001100001000000110100001001100001 :
(key == 11'b00001001000) ? 48'b100000110011001100001101000000110011001100001101 :
(key == 11'b00001001001) ? 48'b100000110010001111000000000000110010001111000000 :
(key == 11'b00001001010) ? 48'b100000110001010001110111000000110001010001110111 :
(key == 11'b00001001011) ? 48'b100000110000010100110011000000110000010100110011 :
(key == 11'b00001001100) ? 48'b100000101111010111110100000000101111010111110100 :
(key == 11'b00001001101) ? 48'b100000101110011010111100000000101110011010111100 :
(key == 11'b00001001110) ? 48'b100000101101011110001001000000101101011110001001 :
(key == 11'b00001001111) ? 48'b100000101100100001011011000000101100100001011011 :
(key == 11'b00001010000) ? 48'b100000101011100100110010000000101011100100110010 :
(key == 11'b00001010001) ? 48'b100000101010101000001110000000101010101000001110 :
(key == 11'b00001010010) ? 48'b100000101001101011110000000000101001101011110000 :
(key == 11'b00001010011) ? 48'b100000101000101111010111000000101000101111010111 :
(key == 11'b00001010100) ? 48'b100000100111110011000011000000100111110011000011 :
(key == 11'b00001010101) ? 48'b100000100110110110110100000000100110110110110100 :
(key == 11'b00001010110) ? 48'b100000100101111010101010000000100101111010101010 :
(key == 11'b00001010111) ? 48'b100000100100111110100111000000100100111110100111 :
(key == 11'b00001011000) ? 48'b100000100100000010101000000000100100000010101000 :
(key == 11'b00001011001) ? 48'b100000100011000110101101000000100011000110101101 :
(key == 11'b00001011010) ? 48'b100000100010001010111000000000100010001010111000 :
(key == 11'b00001011011) ? 48'b100000100001001111001001000000100001001111001001 :
(key == 11'b00001011100) ? 48'b100000100000010011011110000000100000010011011110 :
(key == 11'b00001011101) ? 48'b100000011111010111111001000000011111010111111001 :
(key == 11'b00001011110) ? 48'b100000011110011100011001000000011110011100011001 :
(key == 11'b00001011111) ? 48'b100000011101100000111110000000011101100000111110 :
(key == 11'b00001100000) ? 48'b100000011100100101101000000000011100100101101000 :
(key == 11'b00001100001) ? 48'b100000011011101010010111000000011011101010010111 :
(key == 11'b00001100010) ? 48'b100000011010101111001011000000011010101111001011 :
(key == 11'b00001100011) ? 48'b100000011001110100000100000000011001110100000100 :
(key == 11'b00001100100) ? 48'b100000011000111001000010000000011000111001000010 :
(key == 11'b00001100101) ? 48'b100000010111111110000110000000010111111110000110 :
(key == 11'b00001100110) ? 48'b100000010111000011001110000000010111000011001110 :
(key == 11'b00001100111) ? 48'b100000010110001000011011000000010110001000011011 :
(key == 11'b00001101000) ? 48'b100000010101001101101101000000010101001101101101 :
(key == 11'b00001101001) ? 48'b100000010100010011000101000000010100010011000101 :
(key == 11'b00001101010) ? 48'b100000010011011000100001000000010011011000100001 :
(key == 11'b00001101011) ? 48'b100000010010011110000010000000010010011110000010 :
(key == 11'b00001101100) ? 48'b100000010001100011101000000000010001100011101000 :
(key == 11'b00001101101) ? 48'b100000010000101001010100000000010000101001010100 :
(key == 11'b00001101110) ? 48'b100000001111101111000100000000001111101111000100 :
(key == 11'b00001101111) ? 48'b100000001110110100111000000000001110110100111000 :
(key == 11'b00001110000) ? 48'b100000001101111010110100000000001101111010110100 :
(key == 11'b00001110001) ? 48'b100000001101000000110010000000001101000000110010 :
(key == 11'b00001110010) ? 48'b100000001100000110110101000000001100000110110101 :
(key == 11'b00001110011) ? 48'b100000001011001100111110000000001011001100111110 :
(key == 11'b00001110100) ? 48'b100000001010010011001100000000001010010011001100 :
(key == 11'b00001110101) ? 48'b100000001001011001011101000000001001011001011101 :
(key == 11'b00001110110) ? 48'b100000001000011111110100000000001000011111110100 :
(key == 11'b00001110111) ? 48'b100000000111100110010001000000000111100110010001 :
(key == 11'b00001111000) ? 48'b100000000110101100110001000000000110101100110001 :
(key == 11'b00001111001) ? 48'b100000000101110011010111000000000101110011010111 :
(key == 11'b00001111010) ? 48'b100000000100111010000001000000000100111010000001 :
(key == 11'b00001111011) ? 48'b100000000100000000110001000000000100000000110001 :
(key == 11'b00001111100) ? 48'b100000000011000111100110000000000011000111100110 :
(key == 11'b00001111101) ? 48'b100000000010001110011101000000000010001110011101 :
(key == 11'b00001111110) ? 48'b100000000001010101011011000000000001010101011011 :
(key == 11'b00001111111) ? 48'b100000000000011100011110000000000000011100011110 :
(key == 11'b00010000000) ? 48'b011111111111100011100101111111111111000111001011 :
(key == 11'b00010000001) ? 48'b011111111110101010110001011111111101010101100010 :
(key == 11'b00010000010) ? 48'b011111111101110010000001011111111011100100000010 :
(key == 11'b00010000011) ? 48'b011111111100111001010110011111111001110010101100 :
(key == 11'b00010000100) ? 48'b011111111100000000110000111111111000000001100001 :
(key == 11'b00010000101) ? 48'b011111111011001000001111011111110110010000011110 :
(key == 11'b00010000110) ? 48'b011111111010001111110010111111110100011111100101 :
(key == 11'b00010000111) ? 48'b011111111001010111011010011111110010101110110100 :
(key == 11'b00010001000) ? 48'b011111111000011111000111011111110000111110001110 :
(key == 11'b00010001001) ? 48'b011111110111100110111001111111101111001101110011 :
(key == 11'b00010001010) ? 48'b011111110110101110101111011111101101011101011110 :
(key == 11'b00010001011) ? 48'b011111110101110110101001011111101011101101010010 :
(key == 11'b00010001100) ? 48'b011111110100111110101001011111101001111101010010 :
(key == 11'b00010001101) ? 48'b011111110100000110101100011111101000001101011000 :
(key == 11'b00010001110) ? 48'b011111110011001110110100111111100110011101101001 :
(key == 11'b00010001111) ? 48'b011111110010010111000010111111100100101110000101 :
(key == 11'b00010010000) ? 48'b011111110001011111010011111111100010111110100111 :
(key == 11'b00010010001) ? 48'b011111110000100111101010011111100001001111010100 :
(key == 11'b00010010010) ? 48'b011111101111110000000100111111011111100000001001 :
(key == 11'b00010010011) ? 48'b011111101110111000100100111111011101110001001001 :
(key == 11'b00010010100) ? 48'b011111101110000001001000011111011100000010010000 :
(key == 11'b00010010101) ? 48'b011111101101001001110000111111011010010011100001 :
(key == 11'b00010010110) ? 48'b011111101100010010011101011111011000100100111010 :
(key == 11'b00010010111) ? 48'b011111101011011011001111011111010110110110011110 :
(key == 11'b00010011000) ? 48'b011111101010100100000100011111010101001000001000 :
(key == 11'b00010011001) ? 48'b011111101001101100111111011111010011011001111110 :
(key == 11'b00010011010) ? 48'b011111101000110101111110011111010001101011111100 :
(key == 11'b00010011011) ? 48'b011111100111111111000010011111001111111110000100 :
(key == 11'b00010011100) ? 48'b011111100111001000001010111111001110010000010101 :
(key == 11'b00010011101) ? 48'b011111100110010001010111011111001100100010101110 :
(key == 11'b00010011110) ? 48'b011111100101011010100111111111001010110101001111 :
(key == 11'b00010011111) ? 48'b011111100100100011111100011111001001000111111000 :
(key == 11'b00010100000) ? 48'b011111100011101101010110111111000111011010101101 :
(key == 11'b00010100001) ? 48'b011111100010110110110101011111000101101101101010 :
(key == 11'b00010100010) ? 48'b011111100010000000010111011111000100000000101110 :
(key == 11'b00010100011) ? 48'b011111100001001001111110011111000010010011111100 :
(key == 11'b00010100100) ? 48'b011111100000010011101001011111000000100111010010 :
(key == 11'b00010100101) ? 48'b011111011111011101011000111110111110111010110001 :
(key == 11'b00010100110) ? 48'b011111011110100111001100111110111101001110011001 :
(key == 11'b00010100111) ? 48'b011111011101110001000110011110111011100010001100 :
(key == 11'b00010101000) ? 48'b011111011100111011000010011110111001110110000100 :
(key == 11'b00010101001) ? 48'b011111011100000101000011011110111000001010000110 :
(key == 11'b00010101010) ? 48'b011111011011001111001001011110110110011110010010 :
(key == 11'b00010101011) ? 48'b011111011010011001010010111110110100110010100101 :
(key == 11'b00010101100) ? 48'b011111011001100011100001011110110011000111000010 :
(key == 11'b00010101101) ? 48'b011111011000101101110011111110110001011011100111 :
(key == 11'b00010101110) ? 48'b011111010111111000001010011110101111110000010100 :
(key == 11'b00010101111) ? 48'b011111010111000010100101011110101110000101001010 :
(key == 11'b00010110000) ? 48'b011111010110001101000100111110101100011010001001 :
(key == 11'b00010110001) ? 48'b011111010101010111101000111110101010101111010001 :
(key == 11'b00010110010) ? 48'b011111010100100010001111111110101001000100011111 :
(key == 11'b00010110011) ? 48'b011111010011101100111100011110100111011001111000 :
(key == 11'b00010110100) ? 48'b011111010010110111101100111110100101101111011001 :
(key == 11'b00010110101) ? 48'b011111010010000010100001011110100100000101000010 :
(key == 11'b00010110110) ? 48'b011111010001001101011010011110100010011010110100 :
(key == 11'b00010110111) ? 48'b011111010000011000010111111110100000110000101111 :
(key == 11'b00010111000) ? 48'b011111001111100011011001011110011111000110110010 :
(key == 11'b00010111001) ? 48'b011111001110101110011110111110011101011100111101 :
(key == 11'b00010111010) ? 48'b011111001101111001100111011110011011110011001110 :
(key == 11'b00010111011) ? 48'b011111001101000100110101011110011010001001101010 :
(key == 11'b00010111100) ? 48'b011111001100010000001000111110011000100000010001 :
(key == 11'b00010111101) ? 48'b011111001011011011011111011110010110110110111110 :
(key == 11'b00010111110) ? 48'b011111001010100110111001011110010101001101110010 :
(key == 11'b00010111111) ? 48'b011111001001110010010111011110010011100100101110 :
(key == 11'b00011000000) ? 48'b011111001000111101111010011110010001111011110100 :
(key == 11'b00011000001) ? 48'b011111001000001001100001011110010000010011000010 :
(key == 11'b00011000010) ? 48'b011111000111010101001011111110001110101010010111 :
(key == 11'b00011000011) ? 48'b011111000110100000111011011110001101000001110110 :
(key == 11'b00011000100) ? 48'b011111000101101100101110011110001011011001011100 :
(key == 11'b00011000101) ? 48'b011111000100111000100101011110001001110001001010 :
(key == 11'b00011000110) ? 48'b011111000100000100100001011110001000001001000010 :
(key == 11'b00011000111) ? 48'b011111000011010000100000111110000110100001000001 :
(key == 11'b00011001000) ? 48'b011111000010011100100100111110000100111001001001 :
(key == 11'b00011001001) ? 48'b011111000001101000101011111110000011010001010111 :
(key == 11'b00011001010) ? 48'b011111000000110100111000011110000001101001110000 :
(key == 11'b00011001011) ? 48'b011111000000000001000111011110000000000010001110 :
(key == 11'b00011001100) ? 48'b011110111111001101011011111101111110011010110111 :
(key == 11'b00011001101) ? 48'b011110111110011001110011011101111100110011100110 :
(key == 11'b00011001110) ? 48'b011110111101100110001110011101111011001100011100 :
(key == 11'b00011001111) ? 48'b011110111100110010101111011101111001100101011110 :
(key == 11'b00011010000) ? 48'b011110111011111111010011011101110111111110100110 :
(key == 11'b00011010001) ? 48'b011110111011001011111010011101110110010111110100 :
(key == 11'b00011010010) ? 48'b011110111010011000100111011101110100110001001110 :
(key == 11'b00011010011) ? 48'b011110111001100101010110011101110011001010101100 :
(key == 11'b00011010100) ? 48'b011110111000110010001011011101110001100100010110 :
(key == 11'b00011010101) ? 48'b011110110111111111000011011101101111111110000110 :
(key == 11'b00011010110) ? 48'b011110110111001011111110011101101110010111111100 :
(key == 11'b00011010111) ? 48'b011110110110011000111101111101101100110001111011 :
(key == 11'b00011011000) ? 48'b011110110101100110000010011101101011001100000100 :
(key == 11'b00011011001) ? 48'b011110110100110011001001111101101001100110010011 :
(key == 11'b00011011010) ? 48'b011110110100000000010101011101101000000000101010 :
(key == 11'b00011011011) ? 48'b011110110011001101100100011101100110011011001000 :
(key == 11'b00011011100) ? 48'b011110110010011010111000011101100100110101110000 :
(key == 11'b00011011101) ? 48'b011110110001101000001110111101100011010000011101 :
(key == 11'b00011011110) ? 48'b011110110000110101101011011101100001101011010110 :
(key == 11'b00011011111) ? 48'b011110110000000011001010011101100000000110010100 :
(key == 11'b00011100000) ? 48'b011110101111010000101101011101011110100001011010 :
(key == 11'b00011100001) ? 48'b011110101110011110010100011101011100111100101000 :
(key == 11'b00011100010) ? 48'b011110101101101011111110011101011011010111111100 :
(key == 11'b00011100011) ? 48'b011110101100111001101100111101011001110011011001 :
(key == 11'b00011100100) ? 48'b011110101100000111011111111101011000001110111111 :
(key == 11'b00011100101) ? 48'b011110101011010101010110011101010110101010101100 :
(key == 11'b00011100110) ? 48'b011110101010100011010000011101010101000110100000 :
(key == 11'b00011100111) ? 48'b011110101001110001001101111101010011100010011011 :
(key == 11'b00011101000) ? 48'b011110101000111111001111111101010001111110011111 :
(key == 11'b00011101001) ? 48'b011110101000001101010101011101010000011010101010 :
(key == 11'b00011101010) ? 48'b011110100111011011011111011101001110110110111110 :
(key == 11'b00011101011) ? 48'b011110100110101001101011011101001101010011010110 :
(key == 11'b00011101100) ? 48'b011110100101110111111101011101001011101111111010 :
(key == 11'b00011101101) ? 48'b011110100101000110010010011101001010001100100100 :
(key == 11'b00011101110) ? 48'b011110100100010100101010011101001000101001010100 :
(key == 11'b00011101111) ? 48'b011110100011100011000111011101000111000110001110 :
(key == 11'b00011110000) ? 48'b011110100010110001100111011101000101100011001110 :
(key == 11'b00011110001) ? 48'b011110100010000000001011011101000100000000010110 :
(key == 11'b00011110010) ? 48'b011110100001001110110010111101000010011101100101 :
(key == 11'b00011110011) ? 48'b011110100000011101011110111101000000111010111101 :
(key == 11'b00011110100) ? 48'b011110011111101100001101011100111111011000011010 :
(key == 11'b00011110101) ? 48'b011110011110111010111111111100111101110101111111 :
(key == 11'b00011110110) ? 48'b011110011110001001110111011100111100010011101110 :
(key == 11'b00011110111) ? 48'b011110011101011000110000011100111010110001100000 :
(key == 11'b00011111000) ? 48'b011110011100100111101111011100111001001111011110 :
(key == 11'b00011111001) ? 48'b011110011011110110110001011100110111101101100010 :
(key == 11'b00011111010) ? 48'b011110011011000101110101111100110110001011101011 :
(key == 11'b00011111011) ? 48'b011110011010010100111111011100110100101001111110 :
(key == 11'b00011111100) ? 48'b011110011001100100001100011100110011001000011000 :
(key == 11'b00011111101) ? 48'b011110011000110011011100011100110001100110111000 :
(key == 11'b00011111110) ? 48'b011110011000000010101111111100110000000101011111 :
(key == 11'b00011111111) ? 48'b011110010111010010000111011100101110100100001110 :
(key == 11'b00100000000) ? 48'b011110010110100001100010011100101101000011000100 :
(key == 11'b00100000001) ? 48'b011110010101110001000010011100101011100010000100 :
(key == 11'b00100000010) ? 48'b011110010101000000100101011100101010000001001010 :
(key == 11'b00100000011) ? 48'b011110010100010000001011011100101000100000010110 :
(key == 11'b00100000100) ? 48'b011110010011011111110101011100100110111111101010 :
(key == 11'b00100000101) ? 48'b011110010010101111100010011100100101011111000100 :
(key == 11'b00100000110) ? 48'b011110010001111111010011011100100011111110100110 :
(key == 11'b00100000111) ? 48'b011110010001001111001000011100100010011110010000 :
(key == 11'b00100001000) ? 48'b011110010000011111000001011100100000111110000010 :
(key == 11'b00100001001) ? 48'b011110001111101110111100111100011111011101111001 :
(key == 11'b00100001010) ? 48'b011110001110111110111100011100011101111101111000 :
(key == 11'b00100001011) ? 48'b011110001110001110111111011100011100011101111110 :
(key == 11'b00100001100) ? 48'b011110001101011111000101111100011010111110001011 :
(key == 11'b00100001101) ? 48'b011110001100101111001111011100011001011110011110 :
(key == 11'b00100001110) ? 48'b011110001011111111011101111100010111111110111011 :
(key == 11'b00100001111) ? 48'b011110001011001111101111011100010110011111011110 :
(key == 11'b00100010000) ? 48'b011110001010100000000011011100010101000000000110 :
(key == 11'b00100010001) ? 48'b011110001001110000011011011100010011100000110110 :
(key == 11'b00100010010) ? 48'b011110001001000000110111011100010010000001101110 :
(key == 11'b00100010011) ? 48'b011110001000010001010111011100010000100010101110 :
(key == 11'b00100010100) ? 48'b011110000111100001111001011100001111000011110010 :
(key == 11'b00100010101) ? 48'b011110000110110010100000011100001101100101000000 :
(key == 11'b00100010110) ? 48'b011110000110000011001001011100001100000110010010 :
(key == 11'b00100010111) ? 48'b011110000101010011110111011100001010100111101110 :
(key == 11'b00100011000) ? 48'b011110000100100100100111111100001001001001001111 :
(key == 11'b00100011001) ? 48'b011110000011110101011011011100000111101010110110 :
(key == 11'b00100011010) ? 48'b011110000011000110010011111100000110001100100111 :
(key == 11'b00100011011) ? 48'b011110000010010111001111011100000100101110011110 :
(key == 11'b00100011100) ? 48'b011110000001101000001110011100000011010000011100 :
(key == 11'b00100011101) ? 48'b011110000000111001001111011100000001110010011110 :
(key == 11'b00100011110) ? 48'b011110000000001010010101011100000000010100101010 :
(key == 11'b00100011111) ? 48'b011101111111011011011101111011111110110110111011 :
(key == 11'b00100100000) ? 48'b011101111110101100101010011011111101011001010100 :
(key == 11'b00100100001) ? 48'b011101111101111101111010011011111011111011110100 :
(key == 11'b00100100010) ? 48'b011101111101001111001101011011111010011110011010 :
(key == 11'b00100100011) ? 48'b011101111100100000100100011011111001000001001000 :
(key == 11'b00100100100) ? 48'b011101111011110001111110011011110111100011111100 :
(key == 11'b00100100101) ? 48'b011101111011000011011011111011110110000110110111 :
(key == 11'b00100100110) ? 48'b011101111010010100111100011011110100101001111000 :
(key == 11'b00100100111) ? 48'b011101111001100110100000011011110011001101000000 :
(key == 11'b00100101000) ? 48'b011101111000111000001000011011110001110000010000 :
(key == 11'b00100101001) ? 48'b011101111000001001110011011011110000010011100110 :
(key == 11'b00100101010) ? 48'b011101110111011011100010011011101110110111000100 :
(key == 11'b00100101011) ? 48'b011101110110101101010011011011101101011010100110 :
(key == 11'b00100101100) ? 48'b011101110101111111000111011011101011111110001110 :
(key == 11'b00100101101) ? 48'b011101110101010000111111011011101010100001111110 :
(key == 11'b00100101110) ? 48'b011101110100100010111100011011101001000101111000 :
(key == 11'b00100101111) ? 48'b011101110011110100111010111011100111101001110101 :
(key == 11'b00100110000) ? 48'b011101110011000110111101011011100110001101111010 :
(key == 11'b00100110001) ? 48'b011101110010011001000010111011100100110010000101 :
(key == 11'b00100110010) ? 48'b011101110001101011001100011011100011010110011000 :
(key == 11'b00100110011) ? 48'b011101110000111101011001011011100001111010110010 :
(key == 11'b00100110100) ? 48'b011101110000001111101000011011100000011111010000 :
(key == 11'b00100110101) ? 48'b011101101111100001111010011011011111000011110100 :
(key == 11'b00100110110) ? 48'b011101101110110100010001011011011101101000100010 :
(key == 11'b00100110111) ? 48'b011101101110000110101010011011011100001101010100 :
(key == 11'b00100111000) ? 48'b011101101101011001000111111011011010110010001111 :
(key == 11'b00100111001) ? 48'b011101101100101011100111011011011001010111001110 :
(key == 11'b00100111010) ? 48'b011101101011111110001010011011010111111100010100 :
(key == 11'b00100111011) ? 48'b011101101011010000110001011011010110100001100010 :
(key == 11'b00100111100) ? 48'b011101101010100011011011011011010101000110110110 :
(key == 11'b00100111101) ? 48'b011101101001110110000111011011010011101100001110 :
(key == 11'b00100111110) ? 48'b011101101001001000110111111011010010010001101111 :
(key == 11'b00100111111) ? 48'b011101101000011011101011111011010000110111010111 :
(key == 11'b00101000000) ? 48'b011101100111101110100010011011001111011101000100 :
(key == 11'b00101000001) ? 48'b011101100111000001011100011011001110000010111000 :
(key == 11'b00101000010) ? 48'b011101100110010100011001111011001100101000110011 :
(key == 11'b00101000011) ? 48'b011101100101100111011001111011001011001110110011 :
(key == 11'b00101000100) ? 48'b011101100100111010011101011011001001110100111010 :
(key == 11'b00101000101) ? 48'b011101100100001101100100011011001000011011001000 :
(key == 11'b00101000110) ? 48'b011101100011100000101110011011000111000001011100 :
(key == 11'b00101000111) ? 48'b011101100010110011111011011011000101100111110110 :
(key == 11'b00101001000) ? 48'b011101100010000111001011011011000100001110010110 :
(key == 11'b00101001001) ? 48'b011101100001011010011111011011000010110100111110 :
(key == 11'b00101001010) ? 48'b011101100000101101110110011011000001011011101100 :
(key == 11'b00101001011) ? 48'b011101100000000001001111011011000000000010011110 :
(key == 11'b00101001100) ? 48'b011101011111010100101100111010111110101001011001 :
(key == 11'b00101001101) ? 48'b011101011110101000001101011010111101010000011010 :
(key == 11'b00101001110) ? 48'b011101011101111011110000011010111011110111100000 :
(key == 11'b00101001111) ? 48'b011101011101001111010110011010111010011110101100 :
(key == 11'b00101010000) ? 48'b011101011100100011000000011010111001000110000000 :
(key == 11'b00101010001) ? 48'b011101011011110110101101011010110111101101011010 :
(key == 11'b00101010010) ? 48'b011101011011001010011100111010110110010100111001 :
(key == 11'b00101010011) ? 48'b011101011010011110001111111010110100111100011111 :
(key == 11'b00101010100) ? 48'b011101011001110010000101111010110011100100001011 :
(key == 11'b00101010101) ? 48'b011101011001000101111110111010110010001011111101 :
(key == 11'b00101010110) ? 48'b011101011000011001111010111010110000110011110101 :
(key == 11'b00101010111) ? 48'b011101010111101101111011011010101111011011110110 :
(key == 11'b00101011000) ? 48'b011101010111000001111101011010101110000011111010 :
(key == 11'b00101011001) ? 48'b011101010110010110000010011010101100101100000100 :
(key == 11'b00101011010) ? 48'b011101010101101010001011011010101011010100010110 :
(key == 11'b00101011011) ? 48'b011101010100111110010110111010101001111100101101 :
(key == 11'b00101011100) ? 48'b011101010100010010100101011010101000100101001010 :
(key == 11'b00101011101) ? 48'b011101010011100110110111011010100111001101101110 :
(key == 11'b00101011110) ? 48'b011101010010111011001100011010100101110110011000 :
(key == 11'b00101011111) ? 48'b011101010010001111100011111010100100011111000111 :
(key == 11'b00101100000) ? 48'b011101010001100011111111011010100011000111111110 :
(key == 11'b00101100001) ? 48'b011101010000111000011101011010100001110000111010 :
(key == 11'b00101100010) ? 48'b011101010000001100111110011010100000011001111100 :
(key == 11'b00101100011) ? 48'b011101001111100001100011011010011111000011000110 :
(key == 11'b00101100100) ? 48'b011101001110110110001001011010011101101100010010 :
(key == 11'b00101100101) ? 48'b011101001110001010110011011010011100010101100110 :
(key == 11'b00101100110) ? 48'b011101001101011111011111011010011010111110111110 :
(key == 11'b00101100111) ? 48'b011101001100110100010000011010011001101000100000 :
(key == 11'b00101101000) ? 48'b011101001100001001000011011010011000010010000110 :
(key == 11'b00101101001) ? 48'b011101001011011101111001011010010110111011110010 :
(key == 11'b00101101010) ? 48'b011101001010110010110010111010010101100101100101 :
(key == 11'b00101101011) ? 48'b011101001010000111101110011010010100001111011100 :
(key == 11'b00101101100) ? 48'b011101001001011100101101011010010010111001011010 :
(key == 11'b00101101101) ? 48'b011101001000110001101111111010010001100011011111 :
(key == 11'b00101101110) ? 48'b011101001000000110110100011010010000001101101000 :
(key == 11'b00101101111) ? 48'b011101000111011011111100011010001110110111111000 :
(key == 11'b00101110000) ? 48'b011101000110110001000111111010001101100010001111 :
(key == 11'b00101110001) ? 48'b011101000110000110010101011010001100001100101010 :
(key == 11'b00101110010) ? 48'b011101000101011011100110011010001010110111001100 :
(key == 11'b00101110011) ? 48'b011101000100110000111010011010001001100001110100 :
(key == 11'b00101110100) ? 48'b011101000100000110010000011010001000001100100000 :
(key == 11'b00101110101) ? 48'b011101000011011011101001111010000110110111010011 :
(key == 11'b00101110110) ? 48'b011101000010110001000110011010000101100010001100 :
(key == 11'b00101110111) ? 48'b011101000010000110100101011010000100001101001010 :
(key == 11'b00101111000) ? 48'b011101000001011100001000011010000010111000010000 :
(key == 11'b00101111001) ? 48'b011101000000110001101101011010000001100011011010 :
(key == 11'b00101111010) ? 48'b011101000000000111010110011010000000001110101100 :
(key == 11'b00101111011) ? 48'b011100111111011101000000011001111110111010000000 :
(key == 11'b00101111100) ? 48'b011100111110110010101110011001111101100101011100 :
(key == 11'b00101111101) ? 48'b011100111110001000100000011001111100010001000000 :
(key == 11'b00101111110) ? 48'b011100111101011110010011011001111010111100100110 :
(key == 11'b00101111111) ? 48'b011100111100110100001010011001111001101000010100 :
(key == 11'b00110000000) ? 48'b011100111100001010000011011001111000010100000110 :
(key == 11'b00110000001) ? 48'b011100111011011111111111111001110110111111111111 :
(key == 11'b00110000010) ? 48'b011100111010110101111111011001110101101011111110 :
(key == 11'b00110000011) ? 48'b011100111010001100000001011001110100011000000010 :
(key == 11'b00110000100) ? 48'b011100111001100010000101111001110011000100001011 :
(key == 11'b00110000101) ? 48'b011100111000111000001110011001110001110000011100 :
(key == 11'b00110000110) ? 48'b011100111000001110011000011001110000011100110000 :
(key == 11'b00110000111) ? 48'b011100110111100100100110011001101111001001001100 :
(key == 11'b00110001000) ? 48'b011100110110111010110101111001101101110101101011 :
(key == 11'b00110001001) ? 48'b011100110110010001001001011001101100100010010010 :
(key == 11'b00110001010) ? 48'b011100110101100111011111011001101011001110111110 :
(key == 11'b00110001011) ? 48'b011100110100111101110111111001101001111011101111 :
(key == 11'b00110001100) ? 48'b011100110100010100010010111001101000101000100101 :
(key == 11'b00110001101) ? 48'b011100110011101010110001011001100111010101100010 :
(key == 11'b00110001110) ? 48'b011100110011000001010010011001100110000010100100 :
(key == 11'b00110001111) ? 48'b011100110010010111110110011001100100101111101100 :
(key == 11'b00110010000) ? 48'b011100110001101110011101011001100011011100111010 :
(key == 11'b00110010001) ? 48'b011100110001000101000110111001100010001010001101 :
(key == 11'b00110010010) ? 48'b011100110000011011110011011001100000110111100110 :
(key == 11'b00110010011) ? 48'b011100101111110010100011011001011111100101000110 :
(key == 11'b00110010100) ? 48'b011100101111001001010100011001011110010010101000 :
(key == 11'b00110010101) ? 48'b011100101110100000001001011001011101000000010010 :
(key == 11'b00110010110) ? 48'b011100101101110111000000011001011011101110000000 :
(key == 11'b00110010111) ? 48'b011100101101001101111011011001011010011011110110 :
(key == 11'b00110011000) ? 48'b011100101100100100110111111001011001001001101111 :
(key == 11'b00110011001) ? 48'b011100101011111011110110111001010111110111101101 :
(key == 11'b00110011010) ? 48'b011100101011010010111010011001010110100101110100 :
(key == 11'b00110011011) ? 48'b011100101010101001111110011001010101010011111100 :
(key == 11'b00110011100) ? 48'b011100101010000001000110011001010100000010001100 :
(key == 11'b00110011101) ? 48'b011100101001011000010000111001010010110000100001 :
(key == 11'b00110011110) ? 48'b011100101000101111011110111001010001011110111101 :
(key == 11'b00110011111) ? 48'b011100101000000110101110011001010000001101011100 :
(key == 11'b00110100000) ? 48'b011100100111011110000001011001001110111100000010 :
(key == 11'b00110100001) ? 48'b011100100110110101010111011001001101101010101110 :
(key == 11'b00110100010) ? 48'b011100100110001100101110111001001100011001011101 :
(key == 11'b00110100011) ? 48'b011100100101100100001010011001001011001000010100 :
(key == 11'b00110100100) ? 48'b011100100100111011101000011001001001110111010000 :
(key == 11'b00110100101) ? 48'b011100100100010011001000011001001000100110010000 :
(key == 11'b00110100110) ? 48'b011100100011101010101011011001000111010101010110 :
(key == 11'b00110100111) ? 48'b011100100011000010010001011001000110000100100010 :
(key == 11'b00110101000) ? 48'b011100100010011001111001011001000100110011110010 :
(key == 11'b00110101001) ? 48'b011100100001110001100100011001000011100011001000 :
(key == 11'b00110101010) ? 48'b011100100001001001010010011001000010010010100100 :
(key == 11'b00110101011) ? 48'b011100100000100001000001111001000001000010000011 :
(key == 11'b00110101100) ? 48'b011100011111111000110110011000111111110001101100 :
(key == 11'b00110101101) ? 48'b011100011111010000101011011000111110100001010110 :
(key == 11'b00110101110) ? 48'b011100011110101000100011011000111101010001000110 :
(key == 11'b00110101111) ? 48'b011100011110000000011110011000111100000000111100 :
(key == 11'b00110110000) ? 48'b011100011101011000011011011000111010110000110110 :
(key == 11'b00110110001) ? 48'b011100011100110000011100011000111001100000111000 :
(key == 11'b00110110010) ? 48'b011100011100001000011110111000111000010000111101 :
(key == 11'b00110110011) ? 48'b011100011011100000100101011000110111000001001010 :
(key == 11'b00110110100) ? 48'b011100011010111000101100111000110101110001011001 :
(key == 11'b00110110101) ? 48'b011100011010010000110111011000110100100001101110 :
(key == 11'b00110110110) ? 48'b011100011001101001000100011000110011010010001000 :
(key == 11'b00110110111) ? 48'b011100011001000001010100011000110010000010101000 :
(key == 11'b00110111000) ? 48'b011100011000011001100111011000110000110011001110 :
(key == 11'b00110111001) ? 48'b011100010111110001111100111000101111100011111001 :
(key == 11'b00110111010) ? 48'b011100010111001010010100011000101110010100101000 :
(key == 11'b00110111011) ? 48'b011100010110100010101110111000101101000101011101 :
(key == 11'b00110111100) ? 48'b011100010101111011001011011000101011110110010110 :
(key == 11'b00110111101) ? 48'b011100010101010011101011011000101010100111010110 :
(key == 11'b00110111110) ? 48'b011100010100101100001101011000101001011000011010 :
(key == 11'b00110111111) ? 48'b011100010100000100110010011000101000001001100100 :
(key == 11'b00111000000) ? 48'b011100010011011101011001011000100110111010110010 :
(key == 11'b00111000001) ? 48'b011100010010110110000011011000100101101100000110 :
(key == 11'b00111000010) ? 48'b011100010010001110101111011000100100011101011110 :
(key == 11'b00111000011) ? 48'b011100010001100111011111011000100011001110111110 :
(key == 11'b00111000100) ? 48'b011100010001000000010000011000100010000000100000 :
(key == 11'b00111000101) ? 48'b011100010000011001000011011000100000110010000110 :
(key == 11'b00111000110) ? 48'b011100001111110001111010011000011111100011110100 :
(key == 11'b00111000111) ? 48'b011100001111001010110100011000011110010101101000 :
(key == 11'b00111001000) ? 48'b011100001110100011101111011000011101000111011110 :
(key == 11'b00111001001) ? 48'b011100001101111100101101011000011011111001011010 :
(key == 11'b00111001010) ? 48'b011100001101010101101111011000011010101011011110 :
(key == 11'b00111001011) ? 48'b011100001100101110110010011000011001011101100100 :
(key == 11'b00111001100) ? 48'b011100001100000111111000011000011000001111110000 :
(key == 11'b00111001101) ? 48'b011100001011100000111111011000010111000001111110 :
(key == 11'b00111001110) ? 48'b011100001010111010001010011000010101110100010100 :
(key == 11'b00111001111) ? 48'b011100001010010011011000011000010100100110110000 :
(key == 11'b00111010000) ? 48'b011100001001101100101000011000010011011001010000 :
(key == 11'b00111010001) ? 48'b011100001001000101111010011000010010001011110100 :
(key == 11'b00111010010) ? 48'b011100001000011111001111011000010000111110011110 :
(key == 11'b00111010011) ? 48'b011100000111111000100111011000001111110001001110 :
(key == 11'b00111010100) ? 48'b011100000111010001111111111000001110100011111111 :
(key == 11'b00111010101) ? 48'b011100000110101011011100011000001101010110111000 :
(key == 11'b00111010110) ? 48'b011100000110000100111011111000001100001001110111 :
(key == 11'b00111010111) ? 48'b011100000101011110011100111000001010111100111001 :
(key == 11'b00111011000) ? 48'b011100000100111000000000011000001001110000000000 :
(key == 11'b00111011001) ? 48'b011100000100010001100110011000001000100011001100 :
(key == 11'b00111011010) ? 48'b011100000011101011001110111000000111010110011101 :
(key == 11'b00111011011) ? 48'b011100000011000100111010011000000110001001110100 :
(key == 11'b00111011100) ? 48'b011100000010011110100111011000000100111101001110 :
(key == 11'b00111011101) ? 48'b011100000001111000010111011000000011110000101110 :
(key == 11'b00111011110) ? 48'b011100000001010010001001011000000010100100010010 :
(key == 11'b00111011111) ? 48'b011100000000101011111110111000000001010111111101 :
(key == 11'b00111100000) ? 48'b011100000000000101110101011000000000001011101010 :
(key == 11'b00111100001) ? 48'b011011111111011111110000010111111110111111100000 :
(key == 11'b00111100010) ? 48'b011011111110111001101011010111111101110011010110 :
(key == 11'b00111100011) ? 48'b011011111110010011101010010111111100100111010100 :
(key == 11'b00111100100) ? 48'b011011111101101101101011010111111011011011010110 :
(key == 11'b00111100101) ? 48'b011011111101000111101111010111111010001111011110 :
(key == 11'b00111100110) ? 48'b011011111100100001110100110111111001000011101001 :
(key == 11'b00111100111) ? 48'b011011111011111011111100110111110111110111111001 :
(key == 11'b00111101000) ? 48'b011011111011010110000111110111110110101100001111 :
(key == 11'b00111101001) ? 48'b011011111010110000010101010111110101100000101010 :
(key == 11'b00111101010) ? 48'b011011111010001010100011110111110100010101000111 :
(key == 11'b00111101011) ? 48'b011011111001100100110110010111110011001001101100 :
(key == 11'b00111101100) ? 48'b011011111000111111001010010111110001111110010100 :
(key == 11'b00111101101) ? 48'b011011111000011001100000010111110000110011000000 :
(key == 11'b00111101110) ? 48'b011011110111110011111001110111101111100111110011 :
(key == 11'b00111101111) ? 48'b011011110111001110010101010111101110011100101010 :
(key == 11'b00111110000) ? 48'b011011110110101000110010010111101101010001100100 :
(key == 11'b00111110001) ? 48'b011011110110000011010011010111101100000110100110 :
(key == 11'b00111110010) ? 48'b011011110101011101110110010111101010111011101100 :
(key == 11'b00111110011) ? 48'b011011110100111000011010010111101001110000110100 :
(key == 11'b00111110100) ? 48'b011011110100010011000010010111101000100110000100 :
(key == 11'b00111110101) ? 48'b011011110011101101101011010111100111011011010110 :
(key == 11'b00111110110) ? 48'b011011110011001000010111010111100110010000101110 :
(key == 11'b00111110111) ? 48'b011011110010100011000100010111100101000110001000 :
(key == 11'b00111111000) ? 48'b011011110001111101110101010111100011111011101010 :
(key == 11'b00111111001) ? 48'b011011110001011000101000010111100010110001010000 :
(key == 11'b00111111010) ? 48'b011011110000110011011110010111100001100110111100 :
(key == 11'b00111111011) ? 48'b011011110000001110010101010111100000011100101010 :
(key == 11'b00111111100) ? 48'b011011101111101001001111110111011111010010011111 :
(key == 11'b00111111101) ? 48'b011011101111000100001011010111011110001000010110 :
(key == 11'b00111111110) ? 48'b011011101110011111001001010111011100111110010010 :
(key == 11'b00111111111) ? 48'b011011101101111010001011010111011011110100010110 :
(key == 11'b01000000000) ? 48'b011011101101010101001110010111011010101010011100 :
(key == 11'b01000000001) ? 48'b011011101100110000010011010111011001100000100110 :
(key == 11'b01000000010) ? 48'b011011101100001011011011110111011000010110110111 :
(key == 11'b01000000011) ? 48'b011011101011100110100101110111010111001101001011 :
(key == 11'b01000000100) ? 48'b011011101011000001110010010111010110000011100100 :
(key == 11'b01000000101) ? 48'b011011101010011101000000010111010100111010000000 :
(key == 11'b01000000110) ? 48'b011011101001111000010001010111010011110000100010 :
(key == 11'b01000000111) ? 48'b011011101001010011100100010111010010100111001000 :
(key == 11'b01000001000) ? 48'b011011101000101110111010010111010001011101110100 :
(key == 11'b01000001001) ? 48'b011011101000001010010010010111010000010100100100 :
(key == 11'b01000001010) ? 48'b011011100111100101101100010111001111001011011000 :
(key == 11'b01000001011) ? 48'b011011100111000001001000010111001110000010010000 :
(key == 11'b01000001100) ? 48'b011011100110011100100111010111001100111001001110 :
(key == 11'b01000001101) ? 48'b011011100101111000000111110111001011110000001111 :
(key == 11'b01000001110) ? 48'b011011100101010011101011010111001010100111010110 :
(key == 11'b01000001111) ? 48'b011011100100101111010001010111001001011110100010 :
(key == 11'b01000010000) ? 48'b011011100100001010111000010111001000010101110000 :
(key == 11'b01000010001) ? 48'b011011100011100110100010010111000111001101000100 :
(key == 11'b01000010010) ? 48'b011011100011000010001110010111000110000100011100 :
(key == 11'b01000010011) ? 48'b011011100010011101111101010111000100111011111010 :
(key == 11'b01000010100) ? 48'b011011100001111001101101010111000011110011011010 :
(key == 11'b01000010101) ? 48'b011011100001010101100000010111000010101011000000 :
(key == 11'b01000010110) ? 48'b011011100000110001010101010111000001100010101010 :
(key == 11'b01000010111) ? 48'b011011100000001101001101010111000000011010011010 :
(key == 11'b01000011000) ? 48'b011011011111101001000110010110111111010010001100 :
(key == 11'b01000011001) ? 48'b011011011111000101000001110110111110001010000011 :
(key == 11'b01000011010) ? 48'b011011011110100001000000010110111101000010000000 :
(key == 11'b01000011011) ? 48'b011011011101111101000000010110111011111010000000 :
(key == 11'b01000011100) ? 48'b011011011101011001000010010110111010110010000100 :
(key == 11'b01000011101) ? 48'b011011011100110101000110010110111001101010001100 :
(key == 11'b01000011110) ? 48'b011011011100010001001101110110111000100010011011 :
(key == 11'b01000011111) ? 48'b011011011011101101010110110110110111011010101101 :
(key == 11'b01000100000) ? 48'b011011011011001001100010010110110110010011000100 :
(key == 11'b01000100001) ? 48'b011011011010100101101111010110110101001011011110 :
(key == 11'b01000100010) ? 48'b011011011010000001111111010110110100000011111110 :
(key == 11'b01000100011) ? 48'b011011011001011110010000010110110010111100100000 :
(key == 11'b01000100100) ? 48'b011011011000111010100100110110110001110101001001 :
(key == 11'b01000100101) ? 48'b011011011000010110111010010110110000101101110100 :
(key == 11'b01000100110) ? 48'b011011010111110011010011010110101111100110100110 :
(key == 11'b01000100111) ? 48'b011011010111001111101101010110101110011111011010 :
(key == 11'b01000101000) ? 48'b011011010110101100001010010110101101011000010100 :
(key == 11'b01000101001) ? 48'b011011010110001000101000110110101100010001010001 :
(key == 11'b01000101010) ? 48'b011011010101100101001001110110101011001010010011 :
(key == 11'b01000101011) ? 48'b011011010101000001101101010110101010000011011010 :
(key == 11'b01000101100) ? 48'b011011010100011110010001110110101000111100100011 :
(key == 11'b01000101101) ? 48'b011011010011111010111001010110100111110101110010 :
(key == 11'b01000101110) ? 48'b011011010011010111100010110110100110101111000101 :
(key == 11'b01000101111) ? 48'b011011010010110100001111010110100101101000011110 :
(key == 11'b01000110000) ? 48'b011011010010010000111101010110100100100001111010 :
(key == 11'b01000110001) ? 48'b011011010001101101101101010110100011011011011010 :
(key == 11'b01000110010) ? 48'b011011010001001010011111010110100010010100111110 :
(key == 11'b01000110011) ? 48'b011011010000100111010011010110100001001110100110 :
(key == 11'b01000110100) ? 48'b011011010000000100001001010110100000001000010010 :
(key == 11'b01000110101) ? 48'b011011001111100001000001110110011111000010000011 :
(key == 11'b01000110110) ? 48'b011011001110111101111101010110011101111011111010 :
(key == 11'b01000110111) ? 48'b011011001110011010111001110110011100110101110011 :
(key == 11'b01000111000) ? 48'b011011001101110111111000110110011011101111110001 :
(key == 11'b01000111001) ? 48'b011011001101010100111001010110011010101001110010 :
(key == 11'b01000111010) ? 48'b011011001100110001111100110110011001100011111001 :
(key == 11'b01000111011) ? 48'b011011001100001111000001110110011000011110000011 :
(key == 11'b01000111100) ? 48'b011011001011101100001000010110010111011000010000 :
(key == 11'b01000111101) ? 48'b011011001011001001010010010110010110010010100100 :
(key == 11'b01000111110) ? 48'b011011001010100110011110010110010101001100111100 :
(key == 11'b01000111111) ? 48'b011011001010000011101010110110010100000111010101 :
(key == 11'b01001000000) ? 48'b011011001001100000111011010110010011000001110110 :
(key == 11'b01001000001) ? 48'b011011001000111110001100010110010001111100011000 :
(key == 11'b01001000010) ? 48'b011011001000011011100000010110010000110111000000 :
(key == 11'b01001000011) ? 48'b011011000111111000110110010110001111110001101100 :
(key == 11'b01001000100) ? 48'b011011000111010110001110010110001110101100011100 :
(key == 11'b01001000101) ? 48'b011011000110110011101000010110001101100111010000 :
(key == 11'b01001000110) ? 48'b011011000110010001000100010110001100100010001000 :
(key == 11'b01001000111) ? 48'b011011000101101110100010010110001011011101000100 :
(key == 11'b01001001000) ? 48'b011011000101001100000010010110001010011000000100 :
(key == 11'b01001001001) ? 48'b011011000100101001100101010110001001010011001010 :
(key == 11'b01001001010) ? 48'b011011000100000111001000110110001000001110010001 :
(key == 11'b01001001011) ? 48'b011011000011100100101111010110000111001001011110 :
(key == 11'b01001001100) ? 48'b011011000011000010010111110110000110000100101111 :
(key == 11'b01001001101) ? 48'b011011000010100000000010010110000101000000000100 :
(key == 11'b01001001110) ? 48'b011011000001111101101111010110000011111011011110 :
(key == 11'b01001001111) ? 48'b011011000001011011011110010110000010110110111100 :
(key == 11'b01001010000) ? 48'b011011000000111001001101110110000001110010011011 :
(key == 11'b01001010001) ? 48'b011011000000010111000000010110000000101110000000 :
(key == 11'b01001010010) ? 48'b011010111111110100110101010101111111101001101010 :
(key == 11'b01001010011) ? 48'b011010111111010010101100010101111110100101011000 :
(key == 11'b01001010100) ? 48'b011010111110110000100100110101111101100001001001 :
(key == 11'b01001010101) ? 48'b011010111110001110011111110101111100011100111111 :
(key == 11'b01001010110) ? 48'b011010111101101100011100010101111011011000111000 :
(key == 11'b01001010111) ? 48'b011010111101001010011011010101111010010100110110 :
(key == 11'b01001011000) ? 48'b011010111100101000011100010101111001010000111000 :
(key == 11'b01001011001) ? 48'b011010111100000110011110010101111000001100111100 :
(key == 11'b01001011010) ? 48'b011010111011100100100011010101110111001001000110 :
(key == 11'b01001011011) ? 48'b011010111011000010101010010101110110000101010100 :
(key == 11'b01001011100) ? 48'b011010111010100000110010110101110101000001100101 :
(key == 11'b01001011101) ? 48'b011010111001111110111101010101110011111101111010 :
(key == 11'b01001011110) ? 48'b011010111001011101001010010101110010111010010100 :
(key == 11'b01001011111) ? 48'b011010111000111011011001010101110001110110110010 :
(key == 11'b01001100000) ? 48'b011010111000011001101001110101110000110011010011 :
(key == 11'b01001100001) ? 48'b011010110111110111111100010101101111101111111000 :
(key == 11'b01001100010) ? 48'b011010110111010110010000010101101110101100100000 :
(key == 11'b01001100011) ? 48'b011010110110110100100111010101101101101001001110 :
(key == 11'b01001100100) ? 48'b011010110110010011000000010101101100100110000000 :
(key == 11'b01001100101) ? 48'b011010110101110001011010110101101011100010110101 :
(key == 11'b01001100110) ? 48'b011010110101001111110111010101101010011111101110 :
(key == 11'b01001100111) ? 48'b011010110100101110010110010101101001011100101100 :
(key == 11'b01001101000) ? 48'b011010110100001100110110010101101000011001101100 :
(key == 11'b01001101001) ? 48'b011010110011101011011001010101100111010110110010 :
(key == 11'b01001101010) ? 48'b011010110011001001111110010101100110010011111100 :
(key == 11'b01001101011) ? 48'b011010110010101000100100010101100101010001001000 :
(key == 11'b01001101100) ? 48'b011010110010000111001100010101100100001110011000 :
(key == 11'b01001101101) ? 48'b011010110001100101110110010101100011001011101100 :
(key == 11'b01001101110) ? 48'b011010110001000100100010010101100010001001000100 :
(key == 11'b01001101111) ? 48'b011010110000100011010001010101100001000110100010 :
(key == 11'b01001110000) ? 48'b011010110000000010000001010101100000000100000010 :
(key == 11'b01001110001) ? 48'b011010101111100000110011010101011111000001100110 :
(key == 11'b01001110010) ? 48'b011010101110111111100110010101011101111111001100 :
(key == 11'b01001110011) ? 48'b011010101110011110011101010101011100111100111010 :
(key == 11'b01001110100) ? 48'b011010101101111101010101010101011011111010101010 :
(key == 11'b01001110101) ? 48'b011010101101011100001110010101011010111000011100 :
(key == 11'b01001110110) ? 48'b011010101100111011001010010101011001110110010100 :
(key == 11'b01001110111) ? 48'b011010101100011010000111110101011000110100001111 :
(key == 11'b01001111000) ? 48'b011010101011111001000111010101010111110010001110 :
(key == 11'b01001111001) ? 48'b011010101011011000001000010101010110110000010000 :
(key == 11'b01001111010) ? 48'b011010101010110111001100010101010101101110011000 :
(key == 11'b01001111011) ? 48'b011010101010010110010001010101010100101100100010 :
(key == 11'b01001111100) ? 48'b011010101001110101011000010101010011101010110000 :
(key == 11'b01001111101) ? 48'b011010101001010100100001010101010010101001000010 :
(key == 11'b01001111110) ? 48'b011010101000110011101100010101010001100111011000 :
(key == 11'b01001111111) ? 48'b011010101000010010111010010101010000100101110100 :
(key == 11'b01010000000) ? 48'b011010100111110010000111010101001111100100001110 :
(key == 11'b01010000001) ? 48'b011010100111010001011000110101001110100010110001 :
(key == 11'b01010000010) ? 48'b011010100110110000101010110101001101100001010101 :
(key == 11'b01010000011) ? 48'b011010100110001111111111110101001100011111111111 :
(key == 11'b01010000100) ? 48'b011010100101101111010110010101001011011110101100 :
(key == 11'b01010000101) ? 48'b011010100101001110101101010101001010011101011010 :
(key == 11'b01010000110) ? 48'b011010100100101110000111110101001001011100001111 :
(key == 11'b01010000111) ? 48'b011010100100001101100100010101001000011011001000 :
(key == 11'b01010001000) ? 48'b011010100011101101000010010101000111011010000100 :
(key == 11'b01010001001) ? 48'b011010100011001100100001010101000110011001000010 :
(key == 11'b01010001010) ? 48'b011010100010101100000010010101000101011000000100 :
(key == 11'b01010001011) ? 48'b011010100010001011100110010101000100010111001100 :
(key == 11'b01010001100) ? 48'b011010100001101011001011010101000011010110010110 :
(key == 11'b01010001101) ? 48'b011010100001001010110010010101000010010101100100 :
(key == 11'b01010001110) ? 48'b011010100000101010011011110101000001010100110111 :
(key == 11'b01010001111) ? 48'b011010100000001010000110010101000000010100001100 :
(key == 11'b01010010000) ? 48'b011010011111101001110010010100111111010011100100 :
(key == 11'b01010010001) ? 48'b011010011111001001100001010100111110010011000010 :
(key == 11'b01010010010) ? 48'b011010011110101001010001010100111101010010100010 :
(key == 11'b01010010011) ? 48'b011010011110001001000011010100111100010010000110 :
(key == 11'b01010010100) ? 48'b011010011101101000110111010100111011010001101110 :
(key == 11'b01010010101) ? 48'b011010011101001000101101010100111010010001011010 :
(key == 11'b01010010110) ? 48'b011010011100101000100100110100111001010001001001 :
(key == 11'b01010010111) ? 48'b011010011100001000011110010100111000010000111100 :
(key == 11'b01010011000) ? 48'b011010011011101000011001010100110111010000110010 :
(key == 11'b01010011001) ? 48'b011010011011001000010110010100110110010000101100 :
(key == 11'b01010011010) ? 48'b011010011010101000010110010100110101010000101100 :
(key == 11'b01010011011) ? 48'b011010011010001000010110110100110100010000101101 :
(key == 11'b01010011100) ? 48'b011010011001101000011001010100110011010000110010 :
(key == 11'b01010011101) ? 48'b011010011001001000011101110100110010010000111011 :
(key == 11'b01010011110) ? 48'b011010011000101000100011010100110001010001000110 :
(key == 11'b01010011111) ? 48'b011010011000001000101011010100110000010001010110 :
(key == 11'b01010100000) ? 48'b011010010111101000110101010100101111010001101010 :
(key == 11'b01010100001) ? 48'b011010010111001001000001010100101110010010000010 :
(key == 11'b01010100010) ? 48'b011010010110101001001110010100101101010010011100 :
(key == 11'b01010100011) ? 48'b011010010110001001011101010100101100010010111010 :
(key == 11'b01010100100) ? 48'b011010010101101001101110010100101011010011011100 :
(key == 11'b01010100101) ? 48'b011010010101001010000001010100101010010100000010 :
(key == 11'b01010100110) ? 48'b011010010100101010010101110100101001010100101011 :
(key == 11'b01010100111) ? 48'b011010010100001010101100110100101000010101011001 :
(key == 11'b01010101000) ? 48'b011010010011101011000100010100100111010110001000 :
(key == 11'b01010101001) ? 48'b011010010011001011011101110100100110010110111011 :
(key == 11'b01010101010) ? 48'b011010010010101011111010010100100101010111110100 :
(key == 11'b01010101011) ? 48'b011010010010001100010111010100100100011000101110 :
(key == 11'b01010101100) ? 48'b011010010001101100110111010100100011011001101110 :
(key == 11'b01010101101) ? 48'b011010010001001101010111110100100010011010101111 :
(key == 11'b01010101110) ? 48'b011010010000101101111010110100100001011011110101 :
(key == 11'b01010101111) ? 48'b011010010000001110011111010100100000011100111110 :
(key == 11'b01010110000) ? 48'b011010001111101111000101010100011111011110001010 :
(key == 11'b01010110001) ? 48'b011010001111001111101100110100011110011111011001 :
(key == 11'b01010110010) ? 48'b011010001110110000010110010100011101100000101100 :
(key == 11'b01010110011) ? 48'b011010001110010001000010010100011100100010000100 :
(key == 11'b01010110100) ? 48'b011010001101110001110000010100011011100011100000 :
(key == 11'b01010110101) ? 48'b011010001101010010011111010100011010100100111110 :
(key == 11'b01010110110) ? 48'b011010001100110011010000010100011001100110100000 :
(key == 11'b01010110111) ? 48'b011010001100010100000011010100011000101000000110 :
(key == 11'b01010111000) ? 48'b011010001011110100110111010100010111101001101110 :
(key == 11'b01010111001) ? 48'b011010001011010101101101010100010110101011011010 :
(key == 11'b01010111010) ? 48'b011010001010110110100100010100010101101101001000 :
(key == 11'b01010111011) ? 48'b011010001010010111011101110100010100101110111011 :
(key == 11'b01010111100) ? 48'b011010001001111000011001010100010011110000110010 :
(key == 11'b01010111101) ? 48'b011010001001011001010110010100010010110010101100 :
(key == 11'b01010111110) ? 48'b011010001000111010010100110100010001110100101001 :
(key == 11'b01010111111) ? 48'b011010001000011011010101010100010000110110101010 :
(key == 11'b01011000000) ? 48'b011010000111111100011000010100001111111000110000 :
(key == 11'b01011000001) ? 48'b011010000111011101011011010100001110111010110110 :
(key == 11'b01011000010) ? 48'b011010000110111110100000010100001101111101000000 :
(key == 11'b01011000011) ? 48'b011010000110011111101000010100001100111111010000 :
(key == 11'b01011000100) ? 48'b011010000110000000110001010100001100000001100010 :
(key == 11'b01011000101) ? 48'b011010000101100001111100010100001011000011111000 :
(key == 11'b01011000110) ? 48'b011010000101000011001000010100001010000110010000 :
(key == 11'b01011000111) ? 48'b011010000100100100010110010100001001001000101100 :
(key == 11'b01011001000) ? 48'b011010000100000101100110010100001000001011001100 :
(key == 11'b01011001001) ? 48'b011010000011100110110111010100000111001101101110 :
(key == 11'b01011001010) ? 48'b011010000011001000001011010100000110010000010110 :
(key == 11'b01011001011) ? 48'b011010000010101001011111110100000101010010111111 :
(key == 11'b01011001100) ? 48'b011010000010001010110110010100000100010101101100 :
(key == 11'b01011001101) ? 48'b011010000001101100001110110100000011011000011101 :
(key == 11'b01011001110) ? 48'b011010000001001101101001010100000010011011010010 :
(key == 11'b01011001111) ? 48'b011010000000101111000100010100000001011110001000 :
(key == 11'b01011010000) ? 48'b011010000000010000100010010100000000100001000100 :
(key == 11'b01011010001) ? 48'b011001111111110010000001010011111111100100000010 :
(key == 11'b01011010010) ? 48'b011001111111010011100001010011111110100111000010 :
(key == 11'b01011010011) ? 48'b011001111110110101000100010011111101101010001000 :
(key == 11'b01011010100) ? 48'b011001111110010110100111110011111100101101001111 :
(key == 11'b01011010101) ? 48'b011001111101111000001110010011111011110000011100 :
(key == 11'b01011010110) ? 48'b011001111101011001110101010011111010110011101010 :
(key == 11'b01011010111) ? 48'b011001111100111011011110010011111001110110111100 :
(key == 11'b01011011000) ? 48'b011001111100011101001001010011111000111010010010 :
(key == 11'b01011011001) ? 48'b011001111011111110110101110011110111111101101011 :
(key == 11'b01011011010) ? 48'b011001111011100000100100010011110111000001001000 :
(key == 11'b01011011011) ? 48'b011001111011000010010011010011110110000100100110 :
(key == 11'b01011011100) ? 48'b011001111010100100000101010011110101001000001010 :
(key == 11'b01011011101) ? 48'b011001111010000101111000010011110100001011110000 :
(key == 11'b01011011110) ? 48'b011001111001100111101101010011110011001111011010 :
(key == 11'b01011011111) ? 48'b011001111001001001100010010011110010010011000100 :
(key == 11'b01011100000) ? 48'b011001111000101011011011010011110001010110110110 :
(key == 11'b01011100001) ? 48'b011001111000001101010100010011110000011010101000 :
(key == 11'b01011100010) ? 48'b011001110111101111001111110011101111011110011111 :
(key == 11'b01011100011) ? 48'b011001110111010001001100110011101110100010011001 :
(key == 11'b01011100100) ? 48'b011001110110110011001011010011101101100110010110 :
(key == 11'b01011100101) ? 48'b011001110110010101001011010011101100101010010110 :
(key == 11'b01011100110) ? 48'b011001110101110111001100110011101011101110011001 :
(key == 11'b01011100111) ? 48'b011001110101011001010000010011101010110010100000 :
(key == 11'b01011101000) ? 48'b011001110100111011010101110011101001110110101011 :
(key == 11'b01011101001) ? 48'b011001110100011101011011110011101000111010110111 :
(key == 11'b01011101010) ? 48'b011001110011111111100100010011100111111111001000 :
(key == 11'b01011101011) ? 48'b011001110011100001101101110011100111000011011011 :
(key == 11'b01011101100) ? 48'b011001110011000011111001010011100110000111110010 :
(key == 11'b01011101101) ? 48'b011001110010100110000110010011100101001100001100 :
(key == 11'b01011101110) ? 48'b011001110010001000010101010011100100010000101010 :
(key == 11'b01011101111) ? 48'b011001110001101010100110010011100011010101001100 :
(key == 11'b01011110000) ? 48'b011001110001001100110111010011100010011001101110 :
(key == 11'b01011110001) ? 48'b011001110000101111001011010011100001011110010110 :
(key == 11'b01011110010) ? 48'b011001110000010001100000010011100000100011000000 :
(key == 11'b01011110011) ? 48'b011001101111110011110111110011011111100111101111 :
(key == 11'b01011110100) ? 48'b011001101111010110001111110011011110101100011111 :
(key == 11'b01011110101) ? 48'b011001101110111000101001010011011101110001010010 :
(key == 11'b01011110110) ? 48'b011001101110011011000101010011011100110110001010 :
(key == 11'b01011110111) ? 48'b011001101101111101100011010011011011111011000110 :
(key == 11'b01011111000) ? 48'b011001101101100000000001010011011011000000000010 :
(key == 11'b01011111001) ? 48'b011001101101000010100001010011011010000101000010 :
(key == 11'b01011111010) ? 48'b011001101100100101000011010011011001001010000110 :
(key == 11'b01011111011) ? 48'b011001101100000111100111010011011000001111001110 :
(key == 11'b01011111100) ? 48'b011001101011101010001011110011010111010100010111 :
(key == 11'b01011111101) ? 48'b011001101011001100110010010011010110011001100100 :
(key == 11'b01011111110) ? 48'b011001101010101111011010010011010101011110110100 :
(key == 11'b01011111111) ? 48'b011001101010010010000100010011010100100100001000 :
(key == 11'b01100000000) ? 48'b011001101001110100110000010011010011101001100000 :
(key == 11'b01100000001) ? 48'b011001101001010111011101010011010010101110111010 :
(key == 11'b01100000010) ? 48'b011001101000111010001010110011010001110100010101 :
(key == 11'b01100000011) ? 48'b011001101000011100111010110011010000111001110101 :
(key == 11'b01100000100) ? 48'b011001100111111111101101010011001111111111011010 :
(key == 11'b01100000101) ? 48'b011001100111100010100000010011001111000101000000 :
(key == 11'b01100000110) ? 48'b011001100111000101010101010011001110001010101010 :
(key == 11'b01100000111) ? 48'b011001100110101000001011010011001101010000010110 :
(key == 11'b01100001000) ? 48'b011001100110001011000010110011001100010110000101 :
(key == 11'b01100001001) ? 48'b011001100101101101111100010011001011011011111000 :
(key == 11'b01100001010) ? 48'b011001100101010000110111110011001010100001101111 :
(key == 11'b01100001011) ? 48'b011001100100110011110011110011001001100111100111 :
(key == 11'b01100001100) ? 48'b011001100100010110110010010011001000101101100100 :
(key == 11'b01100001101) ? 48'b011001100011111001110001010011000111110011100010 :
(key == 11'b01100001110) ? 48'b011001100011011100110011010011000110111001100110 :
(key == 11'b01100001111) ? 48'b011001100010111111110101010011000101111111101010 :
(key == 11'b01100010000) ? 48'b011001100010100010111001010011000101000101110010 :
(key == 11'b01100010001) ? 48'b011001100010000101111111110011000100001011111111 :
(key == 11'b01100010010) ? 48'b011001100001101001000111010011000011010010001110 :
(key == 11'b01100010011) ? 48'b011001100001001100001111010011000010011000011110 :
(key == 11'b01100010100) ? 48'b011001100000101111011010010011000001011110110100 :
(key == 11'b01100010101) ? 48'b011001100000010010100101110011000000100101001011 :
(key == 11'b01100010110) ? 48'b011001011111110101110011010010111111101011100110 :
(key == 11'b01100010111) ? 48'b011001011111011001000001110010111110110010000011 :
(key == 11'b01100011000) ? 48'b011001011110111100010010010010111101111000100100 :
(key == 11'b01100011001) ? 48'b011001011110011111100100010010111100111111001000 :
(key == 11'b01100011010) ? 48'b011001011110000010111000010010111100000101110000 :
(key == 11'b01100011011) ? 48'b011001011101100110001101010010111011001100011010 :
(key == 11'b01100011100) ? 48'b011001011101001001100011010010111010010011000110 :
(key == 11'b01100011101) ? 48'b011001011100101100111011010010111001011001110110 :
(key == 11'b01100011110) ? 48'b011001011100010000010101010010111000100000101010 :
(key == 11'b01100011111) ? 48'b011001011011110011110000010010110111100111100000 :
(key == 11'b01100100000) ? 48'b011001011011010111001101010010110110101110011010 :
(key == 11'b01100100001) ? 48'b011001011010111010101010010010110101110101010100 :
(key == 11'b01100100010) ? 48'b011001011010011110001010010010110100111100010100 :
(key == 11'b01100100011) ? 48'b011001011010000001101011010010110100000011010110 :
(key == 11'b01100100100) ? 48'b011001011001100101001101110010110011001010011011 :
(key == 11'b01100100101) ? 48'b011001011001001000110001010010110010010001100010 :
(key == 11'b01100100110) ? 48'b011001011000101100010111010010110001011000101110 :
(key == 11'b01100100111) ? 48'b011001011000001111111110010010110000011111111100 :
(key == 11'b01100101000) ? 48'b011001010111110011100110010010101111100111001100 :
(key == 11'b01100101001) ? 48'b011001010111010111010001010010101110101110100010 :
(key == 11'b01100101010) ? 48'b011001010110111010111100010010101101110101111000 :
(key == 11'b01100101011) ? 48'b011001010110011110101001010010101100111101010010 :
(key == 11'b01100101100) ? 48'b011001010110000010011000010010101100000100110000 :
(key == 11'b01100101101) ? 48'b011001010101100110000111110010101011001100001111 :
(key == 11'b01100101110) ? 48'b011001010101001001111000010010101010010011110000 :
(key == 11'b01100101111) ? 48'b011001010100101101101011110010101001011011010111 :
(key == 11'b01100110000) ? 48'b011001010100010001100000010010101000100011000000 :
(key == 11'b01100110001) ? 48'b011001010011110101010101110010100111101010101011 :
(key == 11'b01100110010) ? 48'b011001010011011001001101010010100110110010011010 :
(key == 11'b01100110011) ? 48'b011001010010111101000101110010100101111010001011 :
(key == 11'b01100110100) ? 48'b011001010010100001000000010010100101000010000000 :
(key == 11'b01100110101) ? 48'b011001010010000100111011110010100100001001110111 :
(key == 11'b01100110110) ? 48'b011001010001101000111001010010100011010001110010 :
(key == 11'b01100110111) ? 48'b011001010001001100110111110010100010011001101111 :
(key == 11'b01100111000) ? 48'b011001010000110000110111010010100001100001101110 :
(key == 11'b01100111001) ? 48'b011001010000010100111000010010100000101001110000 :
(key == 11'b01100111010) ? 48'b011001001111111000111011010010011111110001110110 :
(key == 11'b01100111011) ? 48'b011001001111011101000000010010011110111010000000 :
(key == 11'b01100111100) ? 48'b011001001111000001000101110010011110000010001011 :
(key == 11'b01100111101) ? 48'b011001001110100101001101010010011101001010011010 :
(key == 11'b01100111110) ? 48'b011001001110001001010110010010011100010010101100 :
(key == 11'b01100111111) ? 48'b011001001101101101100000010010011011011011000000 :
(key == 11'b01101000000) ? 48'b011001001101010001101100010010011010100011011000 :
(key == 11'b01101000001) ? 48'b011001001100110101111001010010011001101011110010 :
(key == 11'b01101000010) ? 48'b011001001100011010000111110010011000110100001111 :
(key == 11'b01101000011) ? 48'b011001001011111110010111010010010111111100101110 :
(key == 11'b01101000100) ? 48'b011001001011100010101000010010010111000101010000 :
(key == 11'b01101000101) ? 48'b011001001011000110111011010010010110001101110110 :
(key == 11'b01101000110) ? 48'b011001001010101011001111010010010101010110011110 :
(key == 11'b01101000111) ? 48'b011001001010001111100101010010010100011111001010 :
(key == 11'b01101001000) ? 48'b011001001001110011111100110010010011100111111001 :
(key == 11'b01101001001) ? 48'b011001001001011000010100010010010010110000101000 :
(key == 11'b01101001010) ? 48'b011001001000111100101110010010010001111001011100 :
(key == 11'b01101001011) ? 48'b011001001000100001001001010010010001000010010010 :
(key == 11'b01101001100) ? 48'b011001001000000101100110110010010000001011001101 :
(key == 11'b01101001101) ? 48'b011001000111101010000101010010001111010100001010 :
(key == 11'b01101001110) ? 48'b011001000111001110100100010010001110011101001000 :
(key == 11'b01101001111) ? 48'b011001000110110011000101010010001101100110001010 :
(key == 11'b01101010000) ? 48'b011001000110010111100111010010001100101111001110 :
(key == 11'b01101010001) ? 48'b011001000101111100001010110010001011111000010101 :
(key == 11'b01101010010) ? 48'b011001000101100000110000010010001011000001100000 :
(key == 11'b01101010011) ? 48'b011001000101000101010111010010001010001010101110 :
(key == 11'b01101010100) ? 48'b011001000100101001111111010010001001010011111110 :
(key == 11'b01101010101) ? 48'b011001000100001110101000010010001000011101010000 :
(key == 11'b01101010110) ? 48'b011001000011110011010010110010000111100110100101 :
(key == 11'b01101010111) ? 48'b011001000011010111111111010010000110101111111110 :
(key == 11'b01101011000) ? 48'b011001000010111100101100010010000101111001011000 :
(key == 11'b01101011001) ? 48'b011001000010100001011100010010000101000010111000 :
(key == 11'b01101011010) ? 48'b011001000010000110001100010010000100001100011000 :
(key == 11'b01101011011) ? 48'b011001000001101010111110010010000011010101111100 :
(key == 11'b01101011100) ? 48'b011001000001001111110001010010000010011111100010 :
(key == 11'b01101011101) ? 48'b011001000000110100100101010010000001101001001010 :
(key == 11'b01101011110) ? 48'b011001000000011001011011010010000000110010110110 :
(key == 11'b01101011111) ? 48'b011000111111111110010010010001111111111100100100 :
(key == 11'b01101100000) ? 48'b011000111111100011001011110001111111000110010111 :
(key == 11'b01101100001) ? 48'b011000111111001000000101110001111110010000001011 :
(key == 11'b01101100010) ? 48'b011000111110101101000001010001111101011010000010 :
(key == 11'b01101100011) ? 48'b011000111110010001111101010001111100100011111010 :
(key == 11'b01101100100) ? 48'b011000111101110110111100010001111011101101111000 :
(key == 11'b01101100101) ? 48'b011000111101011011111011010001111010110111110110 :
(key == 11'b01101100110) ? 48'b011000111101000000111100110001111010000001111001 :
(key == 11'b01101100111) ? 48'b011000111100100101111111010001111001001011111110 :
(key == 11'b01101101000) ? 48'b011000111100001011000010110001111000010110000101 :
(key == 11'b01101101001) ? 48'b011000111011110000001000010001110111100000010000 :
(key == 11'b01101101010) ? 48'b011000111011010101001110010001110110101010011100 :
(key == 11'b01101101011) ? 48'b011000111010111010010100110001110101110100101001 :
(key == 11'b01101101100) ? 48'b011000111010011111011110010001110100111110111100 :
(key == 11'b01101101101) ? 48'b011000111010000100101001010001110100001001010010 :
(key == 11'b01101101110) ? 48'b011000111001101001110101010001110011010011101010 :
(key == 11'b01101101111) ? 48'b011000111001001111000010010001110010011110000100 :
(key == 11'b01101110000) ? 48'b011000111000110100010000010001110001101000100000 :
(key == 11'b01101110001) ? 48'b011000111000011001100000010001110000110011000000 :
(key == 11'b01101110010) ? 48'b011000110111111110110001110001101111111101100011 :
(key == 11'b01101110011) ? 48'b011000110111100100000011110001101111001000000111 :
(key == 11'b01101110100) ? 48'b011000110111001001011000010001101110010010110000 :
(key == 11'b01101110101) ? 48'b011000110110101110101101010001101101011101011010 :
(key == 11'b01101110110) ? 48'b011000110110010100000011010001101100101000000110 :
(key == 11'b01101110111) ? 48'b011000110101111001011011010001101011110010110110 :
(key == 11'b01101111000) ? 48'b011000110101011110110101010001101010111101101010 :
(key == 11'b01101111001) ? 48'b011000110101000100001111010001101010001000011110 :
(key == 11'b01101111010) ? 48'b011000110100101001101011010001101001010011010110 :
(key == 11'b01101111011) ? 48'b011000110100001111001000010001101000011110010000 :
(key == 11'b01101111100) ? 48'b011000110011110100100111010001100111101001001110 :
(key == 11'b01101111101) ? 48'b011000110011011010000111010001100110110100001110 :
(key == 11'b01101111110) ? 48'b011000110010111111101000010001100101111111010000 :
(key == 11'b01101111111) ? 48'b011000110010100101001010110001100101001010010101 :
(key == 11'b01110000000) ? 48'b011000110010001010101110110001100100010101011101 :
(key == 11'b01110000001) ? 48'b011000110001110000010011010001100011100000100110 :
(key == 11'b01110000010) ? 48'b011000110001010101111001110001100010101011110011 :
(key == 11'b01110000011) ? 48'b011000110000111011100001010001100001110111000010 :
(key == 11'b01110000100) ? 48'b011000110000100001001011010001100001000010010110 :
(key == 11'b01110000101) ? 48'b011000110000000110110110010001100000001101101100 :
(key == 11'b01110000110) ? 48'b011000101111101100100001110001011111011001000011 :
(key == 11'b01110000111) ? 48'b011000101111010010001110110001011110100100011101 :
(key == 11'b01110001000) ? 48'b011000101110110111111100010001011101101111111000 :
(key == 11'b01110001001) ? 48'b011000101110011101101011110001011100111011010111 :
(key == 11'b01110001010) ? 48'b011000101110000011011101010001011100000110111010 :
(key == 11'b01110001011) ? 48'b011000101101101001001111010001011011010010011110 :
(key == 11'b01110001100) ? 48'b011000101101001111000011010001011010011110000110 :
(key == 11'b01110001101) ? 48'b011000101100110100111000010001011001101001110000 :
(key == 11'b01110001110) ? 48'b011000101100011010101110010001011000110101011100 :
(key == 11'b01110001111) ? 48'b011000101100000000100110010001011000000001001100 :
(key == 11'b01110010000) ? 48'b011000101011100110011110010001010111001100111100 :
(key == 11'b01110010001) ? 48'b011000101011001100011000110001010110011000110001 :
(key == 11'b01110010010) ? 48'b011000101010110010010100110001010101100100101001 :
(key == 11'b01110010011) ? 48'b011000101010011000010001010001010100110000100010 :
(key == 11'b01110010100) ? 48'b011000101001111110001111010001010011111100011110 :
(key == 11'b01110010101) ? 48'b011000101001100100001110010001010011001000011100 :
(key == 11'b01110010110) ? 48'b011000101001001010001110010001010010010100011100 :
(key == 11'b01110010111) ? 48'b011000101000110000010000010001010001100000100000 :
(key == 11'b01110011000) ? 48'b011000101000010110010011010001010000101100100110 :
(key == 11'b01110011001) ? 48'b011000100111111100010111010001001111111000101110 :
(key == 11'b01110011010) ? 48'b011000100111100010011110010001001111000100111100 :
(key == 11'b01110011011) ? 48'b011000100111001000100100010001001110010001001000 :
(key == 11'b01110011100) ? 48'b011000100110101110101100010001001101011101011000 :
(key == 11'b01110011101) ? 48'b011000100110010100110110110001001100101001101101 :
(key == 11'b01110011110) ? 48'b011000100101111011000001010001001011110110000010 :
(key == 11'b01110011111) ? 48'b011000100101100001001101010001001011000010011010 :
(key == 11'b01110100000) ? 48'b011000100101000111011010110001001010001110110101 :
(key == 11'b01110100001) ? 48'b011000100100101101101000110001001001011011010001 :
(key == 11'b01110100010) ? 48'b011000100100010011111001010001001000100111110010 :
(key == 11'b01110100011) ? 48'b011000100011111010001010010001000111110100010100 :
(key == 11'b01110100100) ? 48'b011000100011100000011100010001000111000000111000 :
(key == 11'b01110100101) ? 48'b011000100011000110101111110001000110001101011111 :
(key == 11'b01110100110) ? 48'b011000100010101101000100010001000101011010001000 :
(key == 11'b01110100111) ? 48'b011000100010010011011010110001000100100110110101 :
(key == 11'b01110101000) ? 48'b011000100001111001110001110001000011110011100011 :
(key == 11'b01110101001) ? 48'b011000100001100000001011010001000011000000010110 :
(key == 11'b01110101010) ? 48'b011000100001000110100101010001000010001101001010 :
(key == 11'b01110101011) ? 48'b011000100000101101000000010001000001011010000000 :
(key == 11'b01110101100) ? 48'b011000100000010011011100110001000000100110111001 :
(key == 11'b01110101101) ? 48'b011000011111111001111010010000111111110011110100 :
(key == 11'b01110101110) ? 48'b011000011111100000011001010000111111000000110010 :
(key == 11'b01110101111) ? 48'b011000011111000110111001010000111110001101110010 :
(key == 11'b01110110000) ? 48'b011000011110101101011010010000111101011010110100 :
(key == 11'b01110110001) ? 48'b011000011110010011111101010000111100100111111010 :
(key == 11'b01110110010) ? 48'b011000011101111010100001010000111011110101000010 :
(key == 11'b01110110011) ? 48'b011000011101100001000110010000111011000010001100 :
(key == 11'b01110110100) ? 48'b011000011101000111101100010000111010001111011000 :
(key == 11'b01110110101) ? 48'b011000011100101110010100110000111001011100101001 :
(key == 11'b01110110110) ? 48'b011000011100010100111101110000111000101001111011 :
(key == 11'b01110110111) ? 48'b011000011011111011100111010000110111110111001110 :
(key == 11'b01110111000) ? 48'b011000011011100010010010110000110111000100100101 :
(key == 11'b01110111001) ? 48'b011000011011001000111111010000110110010001111110 :
(key == 11'b01110111010) ? 48'b011000011010101111101101010000110101011111011010 :
(key == 11'b01110111011) ? 48'b011000011010010110011011010000110100101100110110 :
(key == 11'b01110111100) ? 48'b011000011001111101001011110000110011111010010111 :
(key == 11'b01110111101) ? 48'b011000011001100011111101110000110011000111111011 :
(key == 11'b01110111110) ? 48'b011000011001001010110000010000110010010101100000 :
(key == 11'b01110111111) ? 48'b011000011000110001100100010000110001100011001000 :
(key == 11'b01111000000) ? 48'b011000011000011000011001010000110000110000110010 :
(key == 11'b01111000001) ? 48'b011000010111111111001110110000101111111110011101 :
(key == 11'b01111000010) ? 48'b011000010111100110000110110000101111001100001101 :
(key == 11'b01111000011) ? 48'b011000010111001100111110110000101110011001111101 :
(key == 11'b01111000100) ? 48'b011000010110110011111001010000101101100111110010 :
(key == 11'b01111000101) ? 48'b011000010110011010110100110000101100110101101001 :
(key == 11'b01111000110) ? 48'b011000010110000001110000010000101100000011100000 :
(key == 11'b01111000111) ? 48'b011000010101101000101101110000101011010001011011 :
(key == 11'b01111001000) ? 48'b011000010101001111101101010000101010011111011010 :
(key == 11'b01111001001) ? 48'b011000010100110110101100110000101001101101011001 :
(key == 11'b01111001010) ? 48'b011000010100011101101101110000101000111011011011 :
(key == 11'b01111001011) ? 48'b011000010100000100110000010000101000001001100000 :
(key == 11'b01111001100) ? 48'b011000010011101011110100010000100111010111101000 :
(key == 11'b01111001101) ? 48'b011000010011010010111001010000100110100101110010 :
(key == 11'b01111001110) ? 48'b011000010010111001111111010000100101110011111110 :
(key == 11'b01111001111) ? 48'b011000010010100001000110010000100101000010001100 :
(key == 11'b01111010000) ? 48'b011000010010001000001110110000100100010000011101 :
(key == 11'b01111010001) ? 48'b011000010001101111011000110000100011011110110001 :
(key == 11'b01111010010) ? 48'b011000010001010110100010110000100010101101000101 :
(key == 11'b01111010011) ? 48'b011000010000111101101111010000100001111011011110 :
(key == 11'b01111010100) ? 48'b011000010000100100111100010000100001001001111000 :
(key == 11'b01111010101) ? 48'b011000010000001100001010010000100000011000010100 :
(key == 11'b01111010110) ? 48'b011000001111110011011001110000011111100110110011 :
(key == 11'b01111010111) ? 48'b011000001111011010101001110000011110110101010011 :
(key == 11'b01111011000) ? 48'b011000001111000001111100110000011110000011111001 :
(key == 11'b01111011001) ? 48'b011000001110101001001111110000011101010010011111 :
(key == 11'b01111011010) ? 48'b011000001110010000100100010000011100100001001000 :
(key == 11'b01111011011) ? 48'b011000001101110111111000110000011011101111110001 :
(key == 11'b01111011100) ? 48'b011000001101011111001111010000011010111110011110 :
(key == 11'b01111011101) ? 48'b011000001101000110100111010000011010001101001110 :
(key == 11'b01111011110) ? 48'b011000001100101110000000010000011001011100000000 :
(key == 11'b01111011111) ? 48'b011000001100010101011010010000011000101010110100 :
(key == 11'b01111100000) ? 48'b011000001011111100110110010000010111111001101100 :
(key == 11'b01111100001) ? 48'b011000001011100100010010010000010111001000100100 :
(key == 11'b01111100010) ? 48'b011000001011001011110000010000010110010111100000 :
(key == 11'b01111100011) ? 48'b011000001010110011001111010000010101100110011110 :
(key == 11'b01111100100) ? 48'b011000001010011010101111010000010100110101011110 :
(key == 11'b01111100101) ? 48'b011000001010000010010000010000010100000100100000 :
(key == 11'b01111100110) ? 48'b011000001001101001110010010000010011010011100100 :
(key == 11'b01111100111) ? 48'b011000001001010001010101010000010010100010101010 :
(key == 11'b01111101000) ? 48'b011000001000111000111001110000010001110001110011 :
(key == 11'b01111101001) ? 48'b011000001000100000011111010000010001000000111110 :
(key == 11'b01111101010) ? 48'b011000001000001000000110110000010000010000001101 :
(key == 11'b01111101011) ? 48'b011000000111101111101110110000001111011111011101 :
(key == 11'b01111101100) ? 48'b011000000111010111011000010000001110101110110000 :
(key == 11'b01111101101) ? 48'b011000000110111111000010010000001101111110000100 :
(key == 11'b01111101110) ? 48'b011000000110100110101110010000001101001101011100 :
(key == 11'b01111101111) ? 48'b011000000110001110011010110000001100011100110101 :
(key == 11'b01111110000) ? 48'b011000000101110110001000110000001011101100010001 :
(key == 11'b01111110001) ? 48'b011000000101011101110111010000001010111011101110 :
(key == 11'b01111110010) ? 48'b011000000101000101100111110000001010001011001111 :
(key == 11'b01111110011) ? 48'b011000000100101101011000110000001001011010110001 :
(key == 11'b01111110100) ? 48'b011000000100010101001011010000001000101010010110 :
(key == 11'b01111110101) ? 48'b011000000011111100111110010000000111111001111100 :
(key == 11'b01111110110) ? 48'b011000000011100100110011010000000111001001100110 :
(key == 11'b01111110111) ? 48'b011000000011001100101001010000000110011001010010 :
(key == 11'b01111111000) ? 48'b011000000010110100100000010000000101101001000000 :
(key == 11'b01111111001) ? 48'b011000000010011100011000010000000100111000110000 :
(key == 11'b01111111010) ? 48'b011000000010000100010001010000000100001000100010 :
(key == 11'b01111111011) ? 48'b011000000001101100001011010000000011011000010110 :
(key == 11'b01111111100) ? 48'b011000000001010100000111110000000010101000001111 :
(key == 11'b01111111101) ? 48'b011000000000111100000100010000000001111000001000 :
(key == 11'b01111111110) ? 48'b011000000000100100000001110000000001001000000011 :
(key == 11'b01111111111) ? 48'b011000000000001100000001010000000000011000000010 :
(key == 11'b10000000000) ? 48'b101111111111010000000010001111111111010000000010 :
(key == 11'b10000000001) ? 48'b101111111101110000001011001111111101110000001011 :
(key == 11'b10000000010) ? 48'b101111111100010000011101001111111100010000011101 :
(key == 11'b10000000011) ? 48'b101111111010110000111000001111111010110000111000 :
(key == 11'b10000000100) ? 48'b101111111001010001011100001111111001010001011100 :
(key == 11'b10000000101) ? 48'b101111110111110010001000001111110111110010001000 :
(key == 11'b10000000110) ? 48'b101111110110010010111110001111110110010010111110 :
(key == 11'b10000000111) ? 48'b101111110100110011111110001111110100110011111110 :
(key == 11'b10000001000) ? 48'b101111110011010101000100001111110011010101000100 :
(key == 11'b10000001001) ? 48'b101111110001110110010101001111110001110110010101 :
(key == 11'b10000001010) ? 48'b101111110000010111101110001111110000010111101110 :
(key == 11'b10000001011) ? 48'b101111101110111001001110001111101110111001001110 :
(key == 11'b10000001100) ? 48'b101111101101011010111010001111101101011010111010 :
(key == 11'b10000001101) ? 48'b101111101011111100101101001111101011111100101101 :
(key == 11'b10000001110) ? 48'b101111101010011110101000001111101010011110101000 :
(key == 11'b10000001111) ? 48'b101111101001000000101100001111101001000000101100 :
(key == 11'b10000010000) ? 48'b101111100111100010111010001111100111100010111010 :
(key == 11'b10000010001) ? 48'b101111100110000101010000001111100110000101010000 :
(key == 11'b10000010010) ? 48'b101111100100100111101111001111100100100111101111 :
(key == 11'b10000010011) ? 48'b101111100011001010010110001111100011001010010110 :
(key == 11'b10000010100) ? 48'b101111100001101101000110001111100001101101000110 :
(key == 11'b10000010101) ? 48'b101111100000001111111110001111100000001111111110 :
(key == 11'b10000010110) ? 48'b101111011110110010111110001111011110110010111110 :
(key == 11'b10000010111) ? 48'b101111011101010110000111001111011101010110000111 :
(key == 11'b10000011000) ? 48'b101111011011111001011001001111011011111001011001 :
(key == 11'b10000011001) ? 48'b101111011010011100110100001111011010011100110100 :
(key == 11'b10000011010) ? 48'b101111011001000000010111001111011001000000010111 :
(key == 11'b10000011011) ? 48'b101111010111100100000010001111010111100100000010 :
(key == 11'b10000011100) ? 48'b101111010110000111110101001111010110000111110101 :
(key == 11'b10000011101) ? 48'b101111010100101011110001001111010100101011110001 :
(key == 11'b10000011110) ? 48'b101111010011001111110110001111010011001111110110 :
(key == 11'b10000011111) ? 48'b101111010001110100000010001111010001110100000010 :
(key == 11'b10000100000) ? 48'b101111010000011000011000001111010000011000011000 :
(key == 11'b10000100001) ? 48'b101111001110111100110101001111001110111100110101 :
(key == 11'b10000100010) ? 48'b101111001101100001011011001111001101100001011011 :
(key == 11'b10000100011) ? 48'b101111001100000110001010001111001100000110001010 :
(key == 11'b10000100100) ? 48'b101111001010101011000000001111001010101011000000 :
(key == 11'b10000100101) ? 48'b101111001001001111111110001111001001001111111110 :
(key == 11'b10000100110) ? 48'b101111000111110101000110001111000111110101000110 :
(key == 11'b10000100111) ? 48'b101111000110011010010100001111000110011010010100 :
(key == 11'b10000101000) ? 48'b101111000100111111101011001111000100111111101011 :
(key == 11'b10000101001) ? 48'b101111000011100101001010001111000011100101001010 :
(key == 11'b10000101010) ? 48'b101111000010001010110010001111000010001010110010 :
(key == 11'b10000101011) ? 48'b101111000000110000100000001111000000110000100000 :
(key == 11'b10000101100) ? 48'b101110111111010110011001001110111111010110011001 :
(key == 11'b10000101101) ? 48'b101110111101111100011001001110111101111100011001 :
(key == 11'b10000101110) ? 48'b101110111100100010100001001110111100100010100001 :
(key == 11'b10000101111) ? 48'b101110111011001000110001001110111011001000110001 :
(key == 11'b10000110000) ? 48'b101110111001101111001001001110111001101111001001 :
(key == 11'b10000110001) ? 48'b101110111000010101101000001110111000010101101000 :
(key == 11'b10000110010) ? 48'b101110110110111100010001001110110110111100010001 :
(key == 11'b10000110011) ? 48'b101110110101100011000001001110110101100011000001 :
(key == 11'b10000110100) ? 48'b101110110100001001111000001110110100001001111000 :
(key == 11'b10000110101) ? 48'b101110110010110000111001001110110010110000111001 :
(key == 11'b10000110110) ? 48'b101110110001011000000001001110110001011000000001 :
(key == 11'b10000110111) ? 48'b101110101111111111010000001110101111111111010000 :
(key == 11'b10000111000) ? 48'b101110101110100110101000001110101110100110101000 :
(key == 11'b10000111001) ? 48'b101110101101001110001000001110101101001110001000 :
(key == 11'b10000111010) ? 48'b101110101011110101101111001110101011110101101111 :
(key == 11'b10000111011) ? 48'b101110101010011101011110001110101010011101011110 :
(key == 11'b10000111100) ? 48'b101110101001000101010100001110101001000101010100 :
(key == 11'b10000111101) ? 48'b101110100111101101010100001110100111101101010100 :
(key == 11'b10000111110) ? 48'b101110100110010101011010001110100110010101011010 :
(key == 11'b10000111111) ? 48'b101110100100111101101001001110100100111101101001 :
(key == 11'b10001000000) ? 48'b101110100011100110000000001110100011100110000000 :
(key == 11'b10001000001) ? 48'b101110100010001110011101001110100010001110011101 :
(key == 11'b10001000010) ? 48'b101110100000110111000010001110100000110111000010 :
(key == 11'b10001000011) ? 48'b101110011111011111110000001110011111011111110000 :
(key == 11'b10001000100) ? 48'b101110011110001000100100001110011110001000100100 :
(key == 11'b10001000101) ? 48'b101110011100110001100000001110011100110001100000 :
(key == 11'b10001000110) ? 48'b101110011011011010100100001110011011011010100100 :
(key == 11'b10001000111) ? 48'b101110011010000011110000001110011010000011110000 :
(key == 11'b10001001000) ? 48'b101110011000101101000100001110011000101101000100 :
(key == 11'b10001001001) ? 48'b101110010111010110011111001110010111010110011111 :
(key == 11'b10001001010) ? 48'b101110010110000000000010001110010110000000000010 :
(key == 11'b10001001011) ? 48'b101110010100101001101011001110010100101001101011 :
(key == 11'b10001001100) ? 48'b101110010011010011011100001110010011010011011100 :
(key == 11'b10001001101) ? 48'b101110010001111101010110001110010001111101010110 :
(key == 11'b10001001110) ? 48'b101110010000100111010111001110010000100111010111 :
(key == 11'b10001001111) ? 48'b101110001111010001011111001110001111010001011111 :
(key == 11'b10001010000) ? 48'b101110001101111011101111001110001101111011101111 :
(key == 11'b10001010001) ? 48'b101110001100100110000110001110001100100110000110 :
(key == 11'b10001010010) ? 48'b101110001011010000100100001110001011010000100100 :
(key == 11'b10001010011) ? 48'b101110001001111011001010001110001001111011001010 :
(key == 11'b10001010100) ? 48'b101110001000100101110111001110001000100101110111 :
(key == 11'b10001010101) ? 48'b101110000111010000101100001110000111010000101100 :
(key == 11'b10001010110) ? 48'b101110000101111011101000001110000101111011101000 :
(key == 11'b10001010111) ? 48'b101110000100100110101011001110000100100110101011 :
(key == 11'b10001011000) ? 48'b101110000011010001110110001110000011010001110110 :
(key == 11'b10001011001) ? 48'b101110000001111101001000001110000001111101001000 :
(key == 11'b10001011010) ? 48'b101110000000101000100000001110000000101000100000 :
(key == 11'b10001011011) ? 48'b101101111111010100000010001101111111010100000010 :
(key == 11'b10001011100) ? 48'b101101111101111111101010001101111101111111101010 :
(key == 11'b10001011101) ? 48'b101101111100101011011000001101111100101011011000 :
(key == 11'b10001011110) ? 48'b101101111011010111001111001101111011010111001111 :
(key == 11'b10001011111) ? 48'b101101111010000011001100001101111010000011001100 :
(key == 11'b10001100000) ? 48'b101101111000101111010001001101111000101111010001 :
(key == 11'b10001100001) ? 48'b101101110111011011011101001101110111011011011101 :
(key == 11'b10001100010) ? 48'b101101110110000111110000001101110110000111110000 :
(key == 11'b10001100011) ? 48'b101101110100110100001011001101110100110100001011 :
(key == 11'b10001100100) ? 48'b101101110011100000101100001101110011100000101100 :
(key == 11'b10001100101) ? 48'b101101110010001101010101001101110010001101010101 :
(key == 11'b10001100110) ? 48'b101101110000111010000100001101110000111010000100 :
(key == 11'b10001100111) ? 48'b101101101111100110111011001101101111100110111011 :
(key == 11'b10001101000) ? 48'b101101101110010011111000001101101110010011111000 :
(key == 11'b10001101001) ? 48'b101101101101000000111110001101101101000000111110 :
(key == 11'b10001101010) ? 48'b101101101011101110001010001101101011101110001010 :
(key == 11'b10001101011) ? 48'b101101101010011011011100001101101010011011011100 :
(key == 11'b10001101100) ? 48'b101101101001001000110110001101101001001000110110 :
(key == 11'b10001101101) ? 48'b101101100111110110011000001101100111110110011000 :
(key == 11'b10001101110) ? 48'b101101100110100100000000001101100110100100000000 :
(key == 11'b10001101111) ? 48'b101101100101010001101110001101100101010001101110 :
(key == 11'b10001110000) ? 48'b101101100011111111100101001101100011111111100101 :
(key == 11'b10001110001) ? 48'b101101100010101101100001001101100010101101100001 :
(key == 11'b10001110010) ? 48'b101101100001011011100100001101100001011011100100 :
(key == 11'b10001110011) ? 48'b101101100000001001110000001101100000001001110000 :
(key == 11'b10001110100) ? 48'b101101011110111000000001001101011110111000000001 :
(key == 11'b10001110101) ? 48'b101101011101100110011000001101011101100110011000 :
(key == 11'b10001110110) ? 48'b101101011100010100111000001101011100010100111000 :
(key == 11'b10001110111) ? 48'b101101011011000011011110001101011011000011011110 :
(key == 11'b10001111000) ? 48'b101101011001110010001010001101011001110010001010 :
(key == 11'b10001111001) ? 48'b101101011000100000111110001101011000100000111110 :
(key == 11'b10001111010) ? 48'b101101010111001111111000001101010111001111111000 :
(key == 11'b10001111011) ? 48'b101101010101111110111010001101010101111110111010 :
(key == 11'b10001111100) ? 48'b101101010100101110000011001101010100101110000011 :
(key == 11'b10001111101) ? 48'b101101010011011101010001001101010011011101010001 :
(key == 11'b10001111110) ? 48'b101101010010001100100111001101010010001100100111 :
(key == 11'b10001111111) ? 48'b101101010000111100000100001101010000111100000100 :
(key == 11'b10010000000) ? 48'b101101001111101011101000001101001111101011101000 :
(key == 11'b10010000001) ? 48'b101101001110011011010000001101001110011011010000 :
(key == 11'b10010000010) ? 48'b101101001101001011000000001101001101001011000000 :
(key == 11'b10010000011) ? 48'b101101001011111010111000001101001011111010111000 :
(key == 11'b10010000100) ? 48'b101101001010101010110101001101001010101010110101 :
(key == 11'b10010000101) ? 48'b101101001001011010111010001101001001011010111010 :
(key == 11'b10010000110) ? 48'b101101001000001011000100001101001000001011000100 :
(key == 11'b10010000111) ? 48'b101101000110111011010110001101000110111011010110 :
(key == 11'b10010001000) ? 48'b101101000101101011101110001101000101101011101110 :
(key == 11'b10010001001) ? 48'b101101000100011100001110001101000100011100001110 :
(key == 11'b10010001010) ? 48'b101101000011001100110010001101000011001100110010 :
(key == 11'b10010001011) ? 48'b101101000001111101011110001101000001111101011110 :
(key == 11'b10010001100) ? 48'b101101000000101110010001001101000000101110010001 :
(key == 11'b10010001101) ? 48'b101100111111011111001001001100111111011111001001 :
(key == 11'b10010001110) ? 48'b101100111110010000001000001100111110010000001000 :
(key == 11'b10010001111) ? 48'b101100111101000001010000001100111101000001010000 :
(key == 11'b10010010000) ? 48'b101100111011110010011011001100111011110010011011 :
(key == 11'b10010010001) ? 48'b101100111010100011101110001100111010100011101110 :
(key == 11'b10010010010) ? 48'b101100111001010101001000001100111001010101001000 :
(key == 11'b10010010011) ? 48'b101100111000000110101000001100111000000110101000 :
(key == 11'b10010010100) ? 48'b101100110110111000001110001100110110111000001110 :
(key == 11'b10010010101) ? 48'b101100110101101001111010001100110101101001111010 :
(key == 11'b10010010110) ? 48'b101100110100011011101101001100110100011011101101 :
(key == 11'b10010010111) ? 48'b101100110011001101100111001100110011001101100111 :
(key == 11'b10010011000) ? 48'b101100110001111111100110001100110001111111100110 :
(key == 11'b10010011001) ? 48'b101100110000110001101100001100110000110001101100 :
(key == 11'b10010011010) ? 48'b101100101111100011111001001100101111100011111001 :
(key == 11'b10010011011) ? 48'b101100101110010110001100001100101110010110001100 :
(key == 11'b10010011100) ? 48'b101100101101001000100110001100101101001000100110 :
(key == 11'b10010011101) ? 48'b101100101011111011000110001100101011111011000110 :
(key == 11'b10010011110) ? 48'b101100101010101101101011001100101010101101101011 :
(key == 11'b10010011111) ? 48'b101100101001100000010110001100101001100000010110 :
(key == 11'b10010100000) ? 48'b101100101000010011001010001100101000010011001010 :
(key == 11'b10010100001) ? 48'b101100100111000110000010001100100111000110000010 :
(key == 11'b10010100010) ? 48'b101100100101111001000001001100100101111001000001 :
(key == 11'b10010100011) ? 48'b101100100100101100000110001100100100101100000110 :
(key == 11'b10010100100) ? 48'b101100100011011111010001001100100011011111010001 :
(key == 11'b10010100101) ? 48'b101100100010010010100010001100100010010010100010 :
(key == 11'b10010100110) ? 48'b101100100001000101111010001100100001000101111010 :
(key == 11'b10010100111) ? 48'b101100011111111001011000001100011111111001011000 :
(key == 11'b10010101000) ? 48'b101100011110101100111100001100011110101100111100 :
(key == 11'b10010101001) ? 48'b101100011101100000100110001100011101100000100110 :
(key == 11'b10010101010) ? 48'b101100011100010100010110001100011100010100010110 :
(key == 11'b10010101011) ? 48'b101100011011001000001100001100011011001000001100 :
(key == 11'b10010101100) ? 48'b101100011001111100001001001100011001111100001001 :
(key == 11'b10010101101) ? 48'b101100011000110000001100001100011000110000001100 :
(key == 11'b10010101110) ? 48'b101100010111100100010100001100010111100100010100 :
(key == 11'b10010101111) ? 48'b101100010110011000100010001100010110011000100010 :
(key == 11'b10010110000) ? 48'b101100010101001100111000001100010101001100111000 :
(key == 11'b10010110001) ? 48'b101100010100000001010011001100010100000001010011 :
(key == 11'b10010110010) ? 48'b101100010010110101110100001100010010110101110100 :
(key == 11'b10010110011) ? 48'b101100010001101010011010001100010001101010011010 :
(key == 11'b10010110100) ? 48'b101100010000011111001000001100010000011111001000 :
(key == 11'b10010110101) ? 48'b101100001111010011111010001100001111010011111010 :
(key == 11'b10010110110) ? 48'b101100001110001000110011001100001110001000110011 :
(key == 11'b10010110111) ? 48'b101100001100111101110011001100001100111101110011 :
(key == 11'b10010111000) ? 48'b101100001011110010111000001100001011110010111000 :
(key == 11'b10010111001) ? 48'b101100001010101000000011001100001010101000000011 :
(key == 11'b10010111010) ? 48'b101100001001011101010010001100001001011101010010 :
(key == 11'b10010111011) ? 48'b101100001000010010101001001100001000010010101001 :
(key == 11'b10010111100) ? 48'b101100000111001000000111001100000111001000000111 :
(key == 11'b10010111101) ? 48'b101100000101111101101010001100000101111101101010 :
(key == 11'b10010111110) ? 48'b101100000100110011010001001100000100110011010001 :
(key == 11'b10010111111) ? 48'b101100000011101000111111001100000011101000111111 :
(key == 11'b10011000000) ? 48'b101100000010011110110100001100000010011110110100 :
(key == 11'b10011000001) ? 48'b101100000001010100101101001100000001010100101101 :
(key == 11'b10011000010) ? 48'b101100000000001010101101001100000000001010101101 :
(key == 11'b10011000011) ? 48'b101011111111000000110100001011111111000000110100 :
(key == 11'b10011000100) ? 48'b101011111101110110111110001011111101110110111110 :
(key == 11'b10011000101) ? 48'b101011111100101101010000001011111100101101010000 :
(key == 11'b10011000110) ? 48'b101011111011100011100110001011111011100011100110 :
(key == 11'b10011000111) ? 48'b101011111010011010000100001011111010011010000100 :
(key == 11'b10011001000) ? 48'b101011111001010000100110001011111001010000100110 :
(key == 11'b10011001001) ? 48'b101011111000000111001110001011111000000111001110 :
(key == 11'b10011001010) ? 48'b101011110110111101111100001011110110111101111100 :
(key == 11'b10011001011) ? 48'b101011110101110100110000001011110101110100110000 :
(key == 11'b10011001100) ? 48'b101011110100101011101010001011110100101011101010 :
(key == 11'b10011001101) ? 48'b101011110011100010101001001011110011100010101001 :
(key == 11'b10011001110) ? 48'b101011110010011001101110001011110010011001101110 :
(key == 11'b10011001111) ? 48'b101011110001010000111001001011110001010000111001 :
(key == 11'b10011010000) ? 48'b101011110000001000001001001011110000001000001001 :
(key == 11'b10011010001) ? 48'b101011101110111111011110001011101110111111011110 :
(key == 11'b10011010010) ? 48'b101011101101110110111010001011101101110110111010 :
(key == 11'b10011010011) ? 48'b101011101100101110011100001011101100101110011100 :
(key == 11'b10011010100) ? 48'b101011101011100110000100001011101011100110000100 :
(key == 11'b10011010101) ? 48'b101011101010011101110000001011101010011101110000 :
(key == 11'b10011010110) ? 48'b101011101001010101100001001011101001010101100001 :
(key == 11'b10011010111) ? 48'b101011101000001101011000001011101000001101011000 :
(key == 11'b10011011000) ? 48'b101011100111000101010110001011100111000101010110 :
(key == 11'b10011011001) ? 48'b101011100101111101011010001011100101111101011010 :
(key == 11'b10011011010) ? 48'b101011100100110101100001001011100100110101100001 :
(key == 11'b10011011011) ? 48'b101011100011101101101110001011100011101101101110 :
(key == 11'b10011011100) ? 48'b101011100010100110000011001011100010100110000011 :
(key == 11'b10011011101) ? 48'b101011100001011110011100001011100001011110011100 :
(key == 11'b10011011110) ? 48'b101011100000010110111011001011100000010110111011 :
(key == 11'b10011011111) ? 48'b101011011111001111011111001011011111001111011111 :
(key == 11'b10011100000) ? 48'b101011011110001000001000001011011110001000001000 :
(key == 11'b10011100001) ? 48'b101011011101000000111000001011011101000000111000 :
(key == 11'b10011100010) ? 48'b101011011011111001101011001011011011111001101011 :
(key == 11'b10011100011) ? 48'b101011011010110010100101001011011010110010100101 :
(key == 11'b10011100100) ? 48'b101011011001101011100101001011011001101011100101 :
(key == 11'b10011100101) ? 48'b101011011000100100101010001011011000100100101010 :
(key == 11'b10011100110) ? 48'b101011010111011101110100001011010111011101110100 :
(key == 11'b10011100111) ? 48'b101011010110010111000100001011010110010111000100 :
(key == 11'b10011101000) ? 48'b101011010101010000011001001011010101010000011001 :
(key == 11'b10011101001) ? 48'b101011010100001001110011001011010100001001110011 :
(key == 11'b10011101010) ? 48'b101011010011000011010011001011010011000011010011 :
(key == 11'b10011101011) ? 48'b101011010001111100111000001011010001111100111000 :
(key == 11'b10011101100) ? 48'b101011010000110110100011001011010000110110100011 :
(key == 11'b10011101101) ? 48'b101011001111110000010010001011001111110000010010 :
(key == 11'b10011101110) ? 48'b101011001110101010001000001011001110101010001000 :
(key == 11'b10011101111) ? 48'b101011001101100100000011001011001101100100000011 :
(key == 11'b10011110000) ? 48'b101011001100011110000100001011001100011110000100 :
(key == 11'b10011110001) ? 48'b101011001011011000001000001011001011011000001000 :
(key == 11'b10011110010) ? 48'b101011001010010010010011001011001010010010010011 :
(key == 11'b10011110011) ? 48'b101011001001001100100011001011001001001100100011 :
(key == 11'b10011110100) ? 48'b101011001000000110111000001011001000000110111000 :
(key == 11'b10011110101) ? 48'b101011000111000001010010001011000111000001010010 :
(key == 11'b10011110110) ? 48'b101011000101111011110010001011000101111011110010 :
(key == 11'b10011110111) ? 48'b101011000100110110010111001011000100110110010111 :
(key == 11'b10011111000) ? 48'b101011000011110001000001001011000011110001000001 :
(key == 11'b10011111001) ? 48'b101011000010101011110000001011000010101011110000 :
(key == 11'b10011111010) ? 48'b101011000001100110100100001011000001100110100100 :
(key == 11'b10011111011) ? 48'b101011000000100001011110001011000000100001011110 :
(key == 11'b10011111100) ? 48'b101010111111011100011110001010111111011100011110 :
(key == 11'b10011111101) ? 48'b101010111110010111100010001010111110010111100010 :
(key == 11'b10011111110) ? 48'b101010111101010010101011001010111101010010101011 :
(key == 11'b10011111111) ? 48'b101010111100001101111010001010111100001101111010 :
(key == 11'b10100000000) ? 48'b101010111011001001001101001010111011001001001101 :
(key == 11'b10100000001) ? 48'b101010111010000100100110001010111010000100100110 :
(key == 11'b10100000010) ? 48'b101010111001000000000100001010111001000000000100 :
(key == 11'b10100000011) ? 48'b101010110111111011101000001010110111111011101000 :
(key == 11'b10100000100) ? 48'b101010110110110111010000001010110110110111010000 :
(key == 11'b10100000101) ? 48'b101010110101110010111100001010110101110010111100 :
(key == 11'b10100000110) ? 48'b101010110100101110110000001010110100101110110000 :
(key == 11'b10100000111) ? 48'b101010110011101010100111001010110011101010100111 :
(key == 11'b10100001000) ? 48'b101010110010100110100100001010110010100110100100 :
(key == 11'b10100001001) ? 48'b101010110001100010100110001010110001100010100110 :
(key == 11'b10100001010) ? 48'b101010110000011110101101001010110000011110101101 :
(key == 11'b10100001011) ? 48'b101010101111011010111000001010101111011010111000 :
(key == 11'b10100001100) ? 48'b101010101110010111001001001010101110010111001001 :
(key == 11'b10100001101) ? 48'b101010101101010011011110001010101101010011011110 :
(key == 11'b10100001110) ? 48'b101010101100001111111010001010101100001111111010 :
(key == 11'b10100001111) ? 48'b101010101011001100011010001010101011001100011010 :
(key == 11'b10100010000) ? 48'b101010101010001000111110001010101010001000111110 :
(key == 11'b10100010001) ? 48'b101010101001000101101000001010101001000101101000 :
(key == 11'b10100010010) ? 48'b101010101000000010010111001010101000000010010111 :
(key == 11'b10100010011) ? 48'b101010100110111111001100001010100110111111001100 :
(key == 11'b10100010100) ? 48'b101010100101111100000100001010100101111100000100 :
(key == 11'b10100010101) ? 48'b101010100100111001000010001010100100111001000010 :
(key == 11'b10100010110) ? 48'b101010100011110110000100001010100011110110000100 :
(key == 11'b10100010111) ? 48'b101010100010110011001100001010100010110011001100 :
(key == 11'b10100011000) ? 48'b101010100001110000011000001010100001110000011000 :
(key == 11'b10100011001) ? 48'b101010100000101101101010001010100000101101101010 :
(key == 11'b10100011010) ? 48'b101010011111101011000000001010011111101011000000 :
(key == 11'b10100011011) ? 48'b101010011110101000011100001010011110101000011100 :
(key == 11'b10100011100) ? 48'b101010011101100101111100001010011101100101111100 :
(key == 11'b10100011101) ? 48'b101010011100100011100000001010011100100011100000 :
(key == 11'b10100011110) ? 48'b101010011011100001001010001010011011100001001010 :
(key == 11'b10100011111) ? 48'b101010011010011110111000001010011010011110111000 :
(key == 11'b10100100000) ? 48'b101010011001011100101100001010011001011100101100 :
(key == 11'b10100100001) ? 48'b101010011000011010100101001010011000011010100101 :
(key == 11'b10100100010) ? 48'b101010010111011000100010001010010111011000100010 :
(key == 11'b10100100011) ? 48'b101010010110010110100100001010010110010110100100 :
(key == 11'b10100100100) ? 48'b101010010101010100101011001010010101010100101011 :
(key == 11'b10100100101) ? 48'b101010010100010010110111001010010100010010110111 :
(key == 11'b10100100110) ? 48'b101010010011010001001000001010010011010001001000 :
(key == 11'b10100100111) ? 48'b101010010010001111011100001010010010001111011100 :
(key == 11'b10100101000) ? 48'b101010010001001101110111001010010001001101110111 :
(key == 11'b10100101001) ? 48'b101010010000001100010110001010010000001100010110 :
(key == 11'b10100101010) ? 48'b101010001111001010111010001010001111001010111010 :
(key == 11'b10100101011) ? 48'b101010001110001001100001001010001110001001100001 :
(key == 11'b10100101100) ? 48'b101010001101001000001110001010001101001000001110 :
(key == 11'b10100101101) ? 48'b101010001100000110111111001010001100000110111111 :
(key == 11'b10100101110) ? 48'b101010001011000101110110001010001011000101110110 :
(key == 11'b10100101111) ? 48'b101010001010000100110001001010001010000100110001 :
(key == 11'b10100110000) ? 48'b101010001001000011110010001010001001000011110010 :
(key == 11'b10100110001) ? 48'b101010001000000010110110001010001000000010110110 :
(key == 11'b10100110010) ? 48'b101010000111000001111111001010000111000001111111 :
(key == 11'b10100110011) ? 48'b101010000110000001001110001010000110000001001110 :
(key == 11'b10100110100) ? 48'b101010000101000000100000001010000101000000100000 :
(key == 11'b10100110101) ? 48'b101010000011111111110111001010000011111111110111 :
(key == 11'b10100110110) ? 48'b101010000010111111010011001010000010111111010011 :
(key == 11'b10100110111) ? 48'b101010000001111110110011001010000001111110110011 :
(key == 11'b10100111000) ? 48'b101010000000111110011001001010000000111110011001 :
(key == 11'b10100111001) ? 48'b101001111111111110000011001001111111111110000011 :
(key == 11'b10100111010) ? 48'b101001111110111101110001001001111110111101110001 :
(key == 11'b10100111011) ? 48'b101001111101111101100100001001111101111101100100 :
(key == 11'b10100111100) ? 48'b101001111100111101011100001001111100111101011100 :
(key == 11'b10100111101) ? 48'b101001111011111101011000001001111011111101011000 :
(key == 11'b10100111110) ? 48'b101001111010111101011000001001111010111101011000 :
(key == 11'b10100111111) ? 48'b101001111001111101011110001001111001111101011110 :
(key == 11'b10101000000) ? 48'b101001111000111101101000001001111000111101101000 :
(key == 11'b10101000001) ? 48'b101001110111111101110110001001110111111101110110 :
(key == 11'b10101000010) ? 48'b101001110110111110001010001001110110111110001010 :
(key == 11'b10101000011) ? 48'b101001110101111110100001001001110101111110100001 :
(key == 11'b10101000100) ? 48'b101001110100111110111101001001110100111110111101 :
(key == 11'b10101000101) ? 48'b101001110011111111011110001001110011111111011110 :
(key == 11'b10101000110) ? 48'b101001110011000000000011001001110011000000000011 :
(key == 11'b10101000111) ? 48'b101001110010000000101101001001110010000000101101 :
(key == 11'b10101001000) ? 48'b101001110001000001011011001001110001000001011011 :
(key == 11'b10101001001) ? 48'b101001110000000010001110001001110000000010001110 :
(key == 11'b10101001010) ? 48'b101001101111000011000101001001101111000011000101 :
(key == 11'b10101001011) ? 48'b101001101110000100000000001001101110000100000000 :
(key == 11'b10101001100) ? 48'b101001101101000101000000001001101101000101000000 :
(key == 11'b10101001101) ? 48'b101001101100000110000101001001101100000110000101 :
(key == 11'b10101001110) ? 48'b101001101011000111001110001001101011000111001110 :
(key == 11'b10101001111) ? 48'b101001101010001000011100001001101010001000011100 :
(key == 11'b10101010000) ? 48'b101001101001001001101110001001101001001001101110 :
(key == 11'b10101010001) ? 48'b101001101000001011000100001001101000001011000100 :
(key == 11'b10101010010) ? 48'b101001100111001100011110001001100111001100011110 :
(key == 11'b10101010011) ? 48'b101001100110001101111101001001100110001101111101 :
(key == 11'b10101010100) ? 48'b101001100101001111100001001001100101001111100001 :
(key == 11'b10101010101) ? 48'b101001100100010001001001001001100100010001001001 :
(key == 11'b10101010110) ? 48'b101001100011010010110101001001100011010010110101 :
(key == 11'b10101010111) ? 48'b101001100010010100100110001001100010010100100110 :
(key == 11'b10101011000) ? 48'b101001100001010110011011001001100001010110011011 :
(key == 11'b10101011001) ? 48'b101001100000011000010100001001100000011000010100 :
(key == 11'b10101011010) ? 48'b101001011111011010010010001001011111011010010010 :
(key == 11'b10101011011) ? 48'b101001011110011100010100001001011110011100010100 :
(key == 11'b10101011100) ? 48'b101001011101011110011010001001011101011110011010 :
(key == 11'b10101011101) ? 48'b101001011100100000100101001001011100100000100101 :
(key == 11'b10101011110) ? 48'b101001011011100010110100001001011011100010110100 :
(key == 11'b10101011111) ? 48'b101001011010100101000111001001011010100101000111 :
(key == 11'b10101100000) ? 48'b101001011001100111100000001001011001100111100000 :
(key == 11'b10101100001) ? 48'b101001011000101001111011001001011000101001111011 :
(key == 11'b10101100010) ? 48'b101001010111101100011100001001010111101100011100 :
(key == 11'b10101100011) ? 48'b101001010110101111000001001001010110101111000001 :
(key == 11'b10101100100) ? 48'b101001010101110001101001001001010101110001101001 :
(key == 11'b10101100101) ? 48'b101001010100110100010110001001010100110100010110 :
(key == 11'b10101100110) ? 48'b101001010011110111000110001001010011110111000110 :
(key == 11'b10101100111) ? 48'b101001010010111001111100001001010010111001111100 :
(key == 11'b10101101000) ? 48'b101001010001111100110110001001010001111100110110 :
(key == 11'b10101101001) ? 48'b101001010000111111110100001001010000111111110100 :
(key == 11'b10101101010) ? 48'b101001010000000010110111001001010000000010110111 :
(key == 11'b10101101011) ? 48'b101001001111000101111101001001001111000101111101 :
(key == 11'b10101101100) ? 48'b101001001110001001001000001001001110001001001000 :
(key == 11'b10101101101) ? 48'b101001001101001100010111001001001101001100010111 :
(key == 11'b10101101110) ? 48'b101001001100001111101010001001001100001111101010 :
(key == 11'b10101101111) ? 48'b101001001011010011000001001001001011010011000001 :
(key == 11'b10101110000) ? 48'b101001001010010110011101001001001010010110011101 :
(key == 11'b10101110001) ? 48'b101001001001011001111101001001001001011001111101 :
(key == 11'b10101110010) ? 48'b101001001000011101100001001001001000011101100001 :
(key == 11'b10101110011) ? 48'b101001000111100001001001001001000111100001001001 :
(key == 11'b10101110100) ? 48'b101001000110100100110100001001000110100100110100 :
(key == 11'b10101110101) ? 48'b101001000101101000100100001001000101101000100100 :
(key == 11'b10101110110) ? 48'b101001000100101100011001001001000100101100011001 :
(key == 11'b10101110111) ? 48'b101001000011110000010010001001000011110000010010 :
(key == 11'b10101111000) ? 48'b101001000010110100001110001001000010110100001110 :
(key == 11'b10101111001) ? 48'b101001000001111000001111001001000001111000001111 :
(key == 11'b10101111010) ? 48'b101001000000111100010100001001000000111100010100 :
(key == 11'b10101111011) ? 48'b101001000000000000011101001001000000000000011101 :
(key == 11'b10101111100) ? 48'b101000111111000100101010001000111111000100101010 :
(key == 11'b10101111101) ? 48'b101000111110001000111100001000111110001000111100 :
(key == 11'b10101111110) ? 48'b101000111101001101010000001000111101001101010000 :
(key == 11'b10101111111) ? 48'b101000111100010001101010001000111100010001101010 :
(key == 11'b10110000000) ? 48'b101000111011010110000111001000111011010110000111 :
(key == 11'b10110000001) ? 48'b101000111010011010101001001000111010011010101001 :
(key == 11'b10110000010) ? 48'b101000111001011111001110001000111001011111001110 :
(key == 11'b10110000011) ? 48'b101000111000100011111000001000111000100011111000 :
(key == 11'b10110000100) ? 48'b101000110111101000100110001000110111101000100110 :
(key == 11'b10110000101) ? 48'b101000110110101101010111001000110110101101010111 :
(key == 11'b10110000110) ? 48'b101000110101110010001100001000110101110010001100 :
(key == 11'b10110000111) ? 48'b101000110100110111000110001000110100110111000110 :
(key == 11'b10110001000) ? 48'b101000110011111100000100001000110011111100000100 :
(key == 11'b10110001001) ? 48'b101000110011000001000110001000110011000001000110 :
(key == 11'b10110001010) ? 48'b101000110010000110001010001000110010000110001010 :
(key == 11'b10110001011) ? 48'b101000110001001011010100001000110001001011010100 :
(key == 11'b10110001100) ? 48'b101000110000010000100001001000110000010000100001 :
(key == 11'b10110001101) ? 48'b101000101111010101110011001000101111010101110011 :
(key == 11'b10110001110) ? 48'b101000101110011011001000001000101110011011001000 :
(key == 11'b10110001111) ? 48'b101000101101100000100010001000101101100000100010 :
(key == 11'b10110010000) ? 48'b101000101100100110000000001000101100100110000000 :
(key == 11'b10110010001) ? 48'b101000101011101011100001001000101011101011100001 :
(key == 11'b10110010010) ? 48'b101000101010110001000110001000101010110001000110 :
(key == 11'b10110010011) ? 48'b101000101001110110110000001000101001110110110000 :
(key == 11'b10110010100) ? 48'b101000101000111100011101001000101000111100011101 :
(key == 11'b10110010101) ? 48'b101000101000000010001110001000101000000010001110 :
(key == 11'b10110010110) ? 48'b101000100111001000000011001000100111001000000011 :
(key == 11'b10110010111) ? 48'b101000100110001101111100001000100110001101111100 :
(key == 11'b10110011000) ? 48'b101000100101010011111000001000100101010011111000 :
(key == 11'b10110011001) ? 48'b101000100100011001111000001000100100011001111000 :
(key == 11'b10110011010) ? 48'b101000100011011111111110001000100011011111111110 :
(key == 11'b10110011011) ? 48'b101000100010100110000110001000100010100110000110 :
(key == 11'b10110011100) ? 48'b101000100001101100010010001000100001101100010010 :
(key == 11'b10110011101) ? 48'b101000100000110010100010001000100000110010100010 :
(key == 11'b10110011110) ? 48'b101000011111111000110110001000011111111000110110 :
(key == 11'b10110011111) ? 48'b101000011110111111001110001000011110111111001110 :
(key == 11'b10110100000) ? 48'b101000011110000101101010001000011110000101101010 :
(key == 11'b10110100001) ? 48'b101000011101001100001001001000011101001100001001 :
(key == 11'b10110100010) ? 48'b101000011100010010101100001000011100010010101100 :
(key == 11'b10110100011) ? 48'b101000011011011001010100001000011011011001010100 :
(key == 11'b10110100100) ? 48'b101000011010011111111111001000011010011111111111 :
(key == 11'b10110100101) ? 48'b101000011001100110101110001000011001100110101110 :
(key == 11'b10110100110) ? 48'b101000011000101101100000001000011000101101100000 :
(key == 11'b10110100111) ? 48'b101000010111110100010111001000010111110100010111 :
(key == 11'b10110101000) ? 48'b101000010110111011010001001000010110111011010001 :
(key == 11'b10110101001) ? 48'b101000010110000010010000001000010110000010010000 :
(key == 11'b10110101010) ? 48'b101000010101001001010000001000010101001001010000 :
(key == 11'b10110101011) ? 48'b101000010100010000010110001000010100010000010110 :
(key == 11'b10110101100) ? 48'b101000010011010111100000001000010011010111100000 :
(key == 11'b10110101101) ? 48'b101000010010011110101100001000010010011110101100 :
(key == 11'b10110101110) ? 48'b101000010001100101111100001000010001100101111100 :
(key == 11'b10110101111) ? 48'b101000010000101101010010001000010000101101010010 :
(key == 11'b10110110000) ? 48'b101000001111110100101010001000001111110100101010 :
(key == 11'b10110110001) ? 48'b101000001110111100000110001000001110111100000110 :
(key == 11'b10110110010) ? 48'b101000001110000011100110001000001110000011100110 :
(key == 11'b10110110011) ? 48'b101000001101001011001010001000001101001011001010 :
(key == 11'b10110110100) ? 48'b101000001100010010110000001000001100010010110000 :
(key == 11'b10110110101) ? 48'b101000001011011010011010001000001011011010011010 :
(key == 11'b10110110110) ? 48'b101000001010100010001001001000001010100010001001 :
(key == 11'b10110110111) ? 48'b101000001001101001111011001000001001101001111011 :
(key == 11'b10110111000) ? 48'b101000001000110001110001001000001000110001110001 :
(key == 11'b10110111001) ? 48'b101000000111111001101011001000000111111001101011 :
(key == 11'b10110111010) ? 48'b101000000111000001101000001000000111000001101000 :
(key == 11'b10110111011) ? 48'b101000000110001001101001001000000110001001101001 :
(key == 11'b10110111100) ? 48'b101000000101010001101110001000000101010001101110 :
(key == 11'b10110111101) ? 48'b101000000100011001110110001000000100011001110110 :
(key == 11'b10110111110) ? 48'b101000000011100010000010001000000011100010000010 :
(key == 11'b10110111111) ? 48'b101000000010101010010001001000000010101010010001 :
(key == 11'b10111000000) ? 48'b101000000001110010100100001000000001110010100100 :
(key == 11'b10111000001) ? 48'b101000000000111010111100001000000000111010111100 :
(key == 11'b10111000010) ? 48'b101000000000000011010110001000000000000011010110 :
(key == 11'b10111000011) ? 48'b100111111111001011110100000111111111001011110100 :
(key == 11'b10111000100) ? 48'b100111111110010100010110000111111110010100010110 :
(key == 11'b10111000101) ? 48'b100111111101011100111010000111111101011100111010 :
(key == 11'b10111000110) ? 48'b100111111100100101100011000111111100100101100011 :
(key == 11'b10111000111) ? 48'b100111111011101110010000000111111011101110010000 :
(key == 11'b10111001000) ? 48'b100111111010110111000000000111111010110111000000 :
(key == 11'b10111001001) ? 48'b100111111001111111110011000111111001111111110011 :
(key == 11'b10111001010) ? 48'b100111111001001000101011000111111001001000101011 :
(key == 11'b10111001011) ? 48'b100111111000010001100110000111111000010001100110 :
(key == 11'b10111001100) ? 48'b100111110111011010100100000111110111011010100100 :
(key == 11'b10111001101) ? 48'b100111110110100011100101000111110110100011100101 :
(key == 11'b10111001110) ? 48'b100111110101101100101010000111110101101100101010 :
(key == 11'b10111001111) ? 48'b100111110100110101110100000111110100110101110100 :
(key == 11'b10111010000) ? 48'b100111110011111111000001000111110011111111000001 :
(key == 11'b10111010001) ? 48'b100111110011001000010001000111110011001000010001 :
(key == 11'b10111010010) ? 48'b100111110010010001100100000111110010010001100100 :
(key == 11'b10111010011) ? 48'b100111110001011010111100000111110001011010111100 :
(key == 11'b10111010100) ? 48'b100111110000100100010110000111110000100100010110 :
(key == 11'b10111010101) ? 48'b100111101111101101110100000111101111101101110100 :
(key == 11'b10111010110) ? 48'b100111101110110111010110000111101110110111010110 :
(key == 11'b10111010111) ? 48'b100111101110000000111011000111101110000000111011 :
(key == 11'b10111011000) ? 48'b100111101101001010100011000111101101001010100011 :
(key == 11'b10111011001) ? 48'b100111101100010100010000000111101100010100010000 :
(key == 11'b10111011010) ? 48'b100111101011011101111111000111101011011101111111 :
(key == 11'b10111011011) ? 48'b100111101010100111110010000111101010100111110010 :
(key == 11'b10111011100) ? 48'b100111101001110001101000000111101001110001101000 :
(key == 11'b10111011101) ? 48'b100111101000111011100010000111101000111011100010 :
(key == 11'b10111011110) ? 48'b100111101000000101100000000111101000000101100000 :
(key == 11'b10111011111) ? 48'b100111100111001111100001000111100111001111100001 :
(key == 11'b10111100000) ? 48'b100111100110011001100101000111100110011001100101 :
(key == 11'b10111100001) ? 48'b100111100101100011101101000111100101100011101101 :
(key == 11'b10111100010) ? 48'b100111100100101101111000000111100100101101111000 :
(key == 11'b10111100011) ? 48'b100111100011111000000110000111100011111000000110 :
(key == 11'b10111100100) ? 48'b100111100011000010011000000111100011000010011000 :
(key == 11'b10111100101) ? 48'b100111100010001100101110000111100010001100101110 :
(key == 11'b10111100110) ? 48'b100111100001010111000111000111100001010111000111 :
(key == 11'b10111100111) ? 48'b100111100000100001100100000111100000100001100100 :
(key == 11'b10111101000) ? 48'b100111011111101100000011000111011111101100000011 :
(key == 11'b10111101001) ? 48'b100111011110110110100111000111011110110110100111 :
(key == 11'b10111101010) ? 48'b100111011110000001001100000111011110000001001100 :
(key == 11'b10111101011) ? 48'b100111011101001011110110000111011101001011110110 :
(key == 11'b10111101100) ? 48'b100111011100010110100100000111011100010110100100 :
(key == 11'b10111101101) ? 48'b100111011011100001010100000111011011100001010100 :
(key == 11'b10111101110) ? 48'b100111011010101100001000000111011010101100001000 :
(key == 11'b10111101111) ? 48'b100111011001110111000000000111011001110111000000 :
(key == 11'b10111110000) ? 48'b100111011001000001111010000111011001000001111010 :
(key == 11'b10111110001) ? 48'b100111011000001100111001000111011000001100111001 :
(key == 11'b10111110010) ? 48'b100111010111010111111010000111010111010111111010 :
(key == 11'b10111110011) ? 48'b100111010110100010111111000111010110100010111111 :
(key == 11'b10111110100) ? 48'b100111010101101110000111000111010101101110000111 :
(key == 11'b10111110101) ? 48'b100111010100111001010010000111010100111001010010 :
(key == 11'b10111110110) ? 48'b100111010100000100100001000111010100000100100001 :
(key == 11'b10111110111) ? 48'b100111010011001111110010000111010011001111110010 :
(key == 11'b10111111000) ? 48'b100111010010011011001000000111010010011011001000 :
(key == 11'b10111111001) ? 48'b100111010001100110100001000111010001100110100001 :
(key == 11'b10111111010) ? 48'b100111010000110001111101000111010000110001111101 :
(key == 11'b10111111011) ? 48'b100111001111111101011100000111001111111101011100 :
(key == 11'b10111111100) ? 48'b100111001111001000111110000111001111001000111110 :
(key == 11'b10111111101) ? 48'b100111001110010100100100000111001110010100100100 :
(key == 11'b10111111110) ? 48'b100111001101100000001101000111001101100000001101 :
(key == 11'b10111111111) ? 48'b100111001100101011111010000111001100101011111010 :
(key == 11'b11000000000) ? 48'b100111001011110111101001000111001011110111101001 :
(key == 11'b11000000001) ? 48'b100111001011000011011100000111001011000011011100 :
(key == 11'b11000000010) ? 48'b100111001010001111010010000111001010001111010010 :
(key == 11'b11000000011) ? 48'b100111001001011011001100000111001001011011001100 :
(key == 11'b11000000100) ? 48'b100111001000100111001000000111001000100111001000 :
(key == 11'b11000000101) ? 48'b100111000111110011001000000111000111110011001000 :
(key == 11'b11000000110) ? 48'b100111000110111111001011000111000110111111001011 :
(key == 11'b11000000111) ? 48'b100111000110001011010010000111000110001011010010 :
(key == 11'b11000001000) ? 48'b100111000101010111011100000111000101010111011100 :
(key == 11'b11000001001) ? 48'b100111000100100011101000000111000100100011101000 :
(key == 11'b11000001010) ? 48'b100111000011101111111000000111000011101111111000 :
(key == 11'b11000001011) ? 48'b100111000010111100001100000111000010111100001100 :
(key == 11'b11000001100) ? 48'b100111000010001000100010000111000010001000100010 :
(key == 11'b11000001101) ? 48'b100111000001010100111011000111000001010100111011 :
(key == 11'b11000001110) ? 48'b100111000000100001011000000111000000100001011000 :
(key == 11'b11000001111) ? 48'b100110111111101101111000000110111111101101111000 :
(key == 11'b11000010000) ? 48'b100110111110111010011100000110111110111010011100 :
(key == 11'b11000010001) ? 48'b100110111110000111000010000110111110000111000010 :
(key == 11'b11000010010) ? 48'b100110111101010011101100000110111101010011101100 :
(key == 11'b11000010011) ? 48'b100110111100100000011000000110111100100000011000 :
(key == 11'b11000010100) ? 48'b100110111011101101001000000110111011101101001000 :
(key == 11'b11000010101) ? 48'b100110111010111001111011000110111010111001111011 :
(key == 11'b11000010110) ? 48'b100110111010000110110010000110111010000110110010 :
(key == 11'b11000010111) ? 48'b100110111001010011101100000110111001010011101100 :
(key == 11'b11000011000) ? 48'b100110111000100000101000000110111000100000101000 :
(key == 11'b11000011001) ? 48'b100110110111101101100111000110110111101101100111 :
(key == 11'b11000011010) ? 48'b100110110110111010101010000110110110111010101010 :
(key == 11'b11000011011) ? 48'b100110110110000111110000000110110110000111110000 :
(key == 11'b11000011100) ? 48'b100110110101010100111001000110110101010100111001 :
(key == 11'b11000011101) ? 48'b100110110100100010000100000110110100100010000100 :
(key == 11'b11000011110) ? 48'b100110110011101111010100000110110011101111010100 :
(key == 11'b11000011111) ? 48'b100110110010111100100111000110110010111100100111 :
(key == 11'b11000100000) ? 48'b100110110010001001111100000110110010001001111100 :
(key == 11'b11000100001) ? 48'b100110110001010111010100000110110001010111010100 :
(key == 11'b11000100010) ? 48'b100110110000100100110000000110110000100100110000 :
(key == 11'b11000100011) ? 48'b100110101111110010001111000110101111110010001111 :
(key == 11'b11000100100) ? 48'b100110101110111111110001000110101110111111110001 :
(key == 11'b11000100101) ? 48'b100110101110001101010110000110101110001101010110 :
(key == 11'b11000100110) ? 48'b100110101101011010111110000110101101011010111110 :
(key == 11'b11000100111) ? 48'b100110101100101000101001000110101100101000101001 :
(key == 11'b11000101000) ? 48'b100110101011110110010110000110101011110110010110 :
(key == 11'b11000101001) ? 48'b100110101011000100001000000110101011000100001000 :
(key == 11'b11000101010) ? 48'b100110101010010001111100000110101010010001111100 :
(key == 11'b11000101011) ? 48'b100110101001011111110100000110101001011111110100 :
(key == 11'b11000101100) ? 48'b100110101000101101101110000110101000101101101110 :
(key == 11'b11000101101) ? 48'b100110100111111011101011000110100111111011101011 :
(key == 11'b11000101110) ? 48'b100110100111001001101100000110100111001001101100 :
(key == 11'b11000101111) ? 48'b100110100110010111110000000110100110010111110000 :
(key == 11'b11000110000) ? 48'b100110100101100101110110000110100101100101110110 :
(key == 11'b11000110001) ? 48'b100110100100110100000000000110100100110100000000 :
(key == 11'b11000110010) ? 48'b100110100100000010001100000110100100000010001100 :
(key == 11'b11000110011) ? 48'b100110100011010000011100000110100011010000011100 :
(key == 11'b11000110100) ? 48'b100110100010011110101110000110100010011110101110 :
(key == 11'b11000110101) ? 48'b100110100001101101000011000110100001101101000011 :
(key == 11'b11000110110) ? 48'b100110100000111011011100000110100000111011011100 :
(key == 11'b11000110111) ? 48'b100110100000001001111000000110100000001001111000 :
(key == 11'b11000111000) ? 48'b100110011111011000010110000110011111011000010110 :
(key == 11'b11000111001) ? 48'b100110011110100110111000000110011110100110111000 :
(key == 11'b11000111010) ? 48'b100110011101110101011100000110011101110101011100 :
(key == 11'b11000111011) ? 48'b100110011101000100000100000110011101000100000100 :
(key == 11'b11000111100) ? 48'b100110011100010010101110000110011100010010101110 :
(key == 11'b11000111101) ? 48'b100110011011100001011100000110011011100001011100 :
(key == 11'b11000111110) ? 48'b100110011010110000001100000110011010110000001100 :
(key == 11'b11000111111) ? 48'b100110011001111110111111000110011001111110111111 :
(key == 11'b11001000000) ? 48'b100110011001001101110110000110011001001101110110 :
(key == 11'b11001000001) ? 48'b100110011000011100101110000110011000011100101110 :
(key == 11'b11001000010) ? 48'b100110010111101011101010000110010111101011101010 :
(key == 11'b11001000011) ? 48'b100110010110111010101010000110010110111010101010 :
(key == 11'b11001000100) ? 48'b100110010110001001101100000110010110001001101100 :
(key == 11'b11001000101) ? 48'b100110010101011000110001000110010101011000110001 :
(key == 11'b11001000110) ? 48'b100110010100100111111001000110010100100111111001 :
(key == 11'b11001000111) ? 48'b100110010011110111000100000110010011110111000100 :
(key == 11'b11001001000) ? 48'b100110010011000110010000000110010011000110010000 :
(key == 11'b11001001001) ? 48'b100110010010010101100010000110010010010101100010 :
(key == 11'b11001001010) ? 48'b100110010001100100110101000110010001100100110101 :
(key == 11'b11001001011) ? 48'b100110010000110100001100000110010000110100001100 :
(key == 11'b11001001100) ? 48'b100110010000000011100110000110010000000011100110 :
(key == 11'b11001001101) ? 48'b100110001111010011000010000110001111010011000010 :
(key == 11'b11001001110) ? 48'b100110001110100010100000000110001110100010100000 :
(key == 11'b11001001111) ? 48'b100110001101110010000011000110001101110010000011 :
(key == 11'b11001010000) ? 48'b100110001101000001101000000110001101000001101000 :
(key == 11'b11001010001) ? 48'b100110001100010001010000000110001100010001010000 :
(key == 11'b11001010010) ? 48'b100110001011100000111010000110001011100000111010 :
(key == 11'b11001010011) ? 48'b100110001010110000101000000110001010110000101000 :
(key == 11'b11001010100) ? 48'b100110001010000000011000000110001010000000011000 :
(key == 11'b11001010101) ? 48'b100110001001010000001100000110001001010000001100 :
(key == 11'b11001010110) ? 48'b100110001000100000000010000110001000100000000010 :
(key == 11'b11001010111) ? 48'b100110000111101111111010000110000111101111111010 :
(key == 11'b11001011000) ? 48'b100110000110111111110110000110000110111111110110 :
(key == 11'b11001011001) ? 48'b100110000110001111110101000110000110001111110101 :
(key == 11'b11001011010) ? 48'b100110000101011111110110000110000101011111110110 :
(key == 11'b11001011011) ? 48'b100110000100101111111010000110000100101111111010 :
(key == 11'b11001011100) ? 48'b100110000100000000000010000110000100000000000010 :
(key == 11'b11001011101) ? 48'b100110000011010000001011000110000011010000001011 :
(key == 11'b11001011110) ? 48'b100110000010100000011000000110000010100000011000 :
(key == 11'b11001011111) ? 48'b100110000001110000100111000110000001110000100111 :
(key == 11'b11001100000) ? 48'b100110000001000000111001000110000001000000111001 :
(key == 11'b11001100001) ? 48'b100110000000010001001110000110000000010001001110 :
(key == 11'b11001100010) ? 48'b100101111111100001100110000101111111100001100110 :
(key == 11'b11001100011) ? 48'b100101111110110010000001000101111110110010000001 :
(key == 11'b11001100100) ? 48'b100101111110000010011111000101111110000010011111 :
(key == 11'b11001100101) ? 48'b100101111101010010111110000101111101010010111110 :
(key == 11'b11001100110) ? 48'b100101111100100011100010000101111100100011100010 :
(key == 11'b11001100111) ? 48'b100101111011110100001000000101111011110100001000 :
(key == 11'b11001101000) ? 48'b100101111011000100110000000101111011000100110000 :
(key == 11'b11001101001) ? 48'b100101111010010101011100000101111010010101011100 :
(key == 11'b11001101010) ? 48'b100101111001100110001010000101111001100110001010 :
(key == 11'b11001101011) ? 48'b100101111000110110111100000101111000110110111100 :
(key == 11'b11001101100) ? 48'b100101111000000111101111000101111000000111101111 :
(key == 11'b11001101101) ? 48'b100101110111011000100101000101110111011000100101 :
(key == 11'b11001101110) ? 48'b100101110110101001011110000101110110101001011110 :
(key == 11'b11001101111) ? 48'b100101110101111010011011000101110101111010011011 :
(key == 11'b11001110000) ? 48'b100101110101001011011010000101110101001011011010 :
(key == 11'b11001110001) ? 48'b100101110100011100011011000101110100011100011011 :
(key == 11'b11001110010) ? 48'b100101110011101101011110000101110011101101011110 :
(key == 11'b11001110011) ? 48'b100101110010111110100110000101110010111110100110 :
(key == 11'b11001110100) ? 48'b100101110010001111110000000101110010001111110000 :
(key == 11'b11001110101) ? 48'b100101110001100000111100000101110001100000111100 :
(key == 11'b11001110110) ? 48'b100101110000110010001010000101110000110010001010 :
(key == 11'b11001110111) ? 48'b100101110000000011011100000101110000000011011100 :
(key == 11'b11001111000) ? 48'b100101101111010100110001000101101111010100110001 :
(key == 11'b11001111001) ? 48'b100101101110100110001000000101101110100110001000 :
(key == 11'b11001111010) ? 48'b100101101101110111100010000101101101110111100010 :
(key == 11'b11001111011) ? 48'b100101101101001000111111000101101101001000111111 :
(key == 11'b11001111100) ? 48'b100101101100011010011110000101101100011010011110 :
(key == 11'b11001111101) ? 48'b100101101011101100000000000101101011101100000000 :
(key == 11'b11001111110) ? 48'b100101101010111101100101000101101010111101100101 :
(key == 11'b11001111111) ? 48'b100101101010001111001100000101101010001111001100 :
(key == 11'b11010000000) ? 48'b100101101001100000110110000101101001100000110110 :
(key == 11'b11010000001) ? 48'b100101101000110010100011000101101000110010100011 :
(key == 11'b11010000010) ? 48'b100101101000000100010010000101101000000100010010 :
(key == 11'b11010000011) ? 48'b100101100111010110000100000101100111010110000100 :
(key == 11'b11010000100) ? 48'b100101100110100111111001000101100110100111111001 :
(key == 11'b11010000101) ? 48'b100101100101111001110000000101100101111001110000 :
(key == 11'b11010000110) ? 48'b100101100101001011101010000101100101001011101010 :
(key == 11'b11010000111) ? 48'b100101100100011101100111000101100100011101100111 :
(key == 11'b11010001000) ? 48'b100101100011101111100110000101100011101111100110 :
(key == 11'b11010001001) ? 48'b100101100011000001101000000101100011000001101000 :
(key == 11'b11010001010) ? 48'b100101100010010011101100000101100010010011101100 :
(key == 11'b11010001011) ? 48'b100101100001100101110011000101100001100101110011 :
(key == 11'b11010001100) ? 48'b100101100000110111111101000101100000110111111101 :
(key == 11'b11010001101) ? 48'b100101100000001010001010000101100000001010001010 :
(key == 11'b11010001110) ? 48'b100101011111011100011010000101011111011100011010 :
(key == 11'b11010001111) ? 48'b100101011110101110101011000101011110101110101011 :
(key == 11'b11010010000) ? 48'b100101011110000000111110000101011110000000111110 :
(key == 11'b11010010001) ? 48'b100101011101010011010110000101011101010011010110 :
(key == 11'b11010010010) ? 48'b100101011100100101101111000101011100100101101111 :
(key == 11'b11010010011) ? 48'b100101011011111000001011000101011011111000001011 :
(key == 11'b11010010100) ? 48'b100101011011001010101010000101011011001010101010 :
(key == 11'b11010010101) ? 48'b100101011010011101001011000101011010011101001011 :
(key == 11'b11010010110) ? 48'b100101011001101111101111000101011001101111101111 :
(key == 11'b11010010111) ? 48'b100101011001000010010110000101011001000010010110 :
(key == 11'b11010011000) ? 48'b100101011000010100111110000101011000010100111110 :
(key == 11'b11010011001) ? 48'b100101010111100111101010000101010111100111101010 :
(key == 11'b11010011010) ? 48'b100101010110111010011001000101010110111010011001 :
(key == 11'b11010011011) ? 48'b100101010110001101001001000101010110001101001001 :
(key == 11'b11010011100) ? 48'b100101010101011111111101000101010101011111111101 :
(key == 11'b11010011101) ? 48'b100101010100110010110010000101010100110010110010 :
(key == 11'b11010011110) ? 48'b100101010100000101101011000101010100000101101011 :
(key == 11'b11010011111) ? 48'b100101010011011000100110000101010011011000100110 :
(key == 11'b11010100000) ? 48'b100101010010101011100011000101010010101011100011 :
(key == 11'b11010100001) ? 48'b100101010001111110100100000101010001111110100100 :
(key == 11'b11010100010) ? 48'b100101010001010001100110000101010001010001100110 :
(key == 11'b11010100011) ? 48'b100101010000100100101011000101010000100100101011 :
(key == 11'b11010100100) ? 48'b100101001111110111110010000101001111110111110010 :
(key == 11'b11010100101) ? 48'b100101001111001010111101000101001111001010111101 :
(key == 11'b11010100110) ? 48'b100101001110011110001010000101001110011110001010 :
(key == 11'b11010100111) ? 48'b100101001101110001011010000101001101110001011010 :
(key == 11'b11010101000) ? 48'b100101001101000100101100000101001101000100101100 :
(key == 11'b11010101001) ? 48'b100101001100010111111111000101001100010111111111 :
(key == 11'b11010101010) ? 48'b100101001011101011010110000101001011101011010110 :
(key == 11'b11010101011) ? 48'b100101001010111110101111000101001010111110101111 :
(key == 11'b11010101100) ? 48'b100101001010010010001100000101001010010010001100 :
(key == 11'b11010101101) ? 48'b100101001001100101101010000101001001100101101010 :
(key == 11'b11010101110) ? 48'b100101001000111001001010000101001000111001001010 :
(key == 11'b11010101111) ? 48'b100101001000001100101110000101001000001100101110 :
(key == 11'b11010110000) ? 48'b100101000111100000010100000101000111100000010100 :
(key == 11'b11010110001) ? 48'b100101000110110011111100000101000110110011111100 :
(key == 11'b11010110010) ? 48'b100101000110000111100110000101000110000111100110 :
(key == 11'b11010110011) ? 48'b100101000101011011010100000101000101011011010100 :
(key == 11'b11010110100) ? 48'b100101000100101111000100000101000100101111000100 :
(key == 11'b11010110101) ? 48'b100101000100000010110110000101000100000010110110 :
(key == 11'b11010110110) ? 48'b100101000011010110101011000101000011010110101011 :
(key == 11'b11010110111) ? 48'b100101000010101010100010000101000010101010100010 :
(key == 11'b11010111000) ? 48'b100101000001111110011100000101000001111110011100 :
(key == 11'b11010111001) ? 48'b100101000001010010011000000101000001010010011000 :
(key == 11'b11010111010) ? 48'b100101000000100110010110000101000000100110010110 :
(key == 11'b11010111011) ? 48'b100100111111111010010111000100111111111010010111 :
(key == 11'b11010111100) ? 48'b100100111111001110011011000100111111001110011011 :
(key == 11'b11010111101) ? 48'b100100111110100010100001000100111110100010100001 :
(key == 11'b11010111110) ? 48'b100100111101110110101001000100111101110110101001 :
(key == 11'b11010111111) ? 48'b100100111101001010110100000100111101001010110100 :
(key == 11'b11011000000) ? 48'b100100111100011111000010000100111100011111000010 :
(key == 11'b11011000001) ? 48'b100100111011110011010010000100111011110011010010 :
(key == 11'b11011000010) ? 48'b100100111011000111100010000100111011000111100010 :
(key == 11'b11011000011) ? 48'b100100111010011011110111000100111010011011110111 :
(key == 11'b11011000100) ? 48'b100100111001110000001110000100111001110000001110 :
(key == 11'b11011000101) ? 48'b100100111001000100101000000100111001000100101000 :
(key == 11'b11011000110) ? 48'b100100111000011001000100000100111000011001000100 :
(key == 11'b11011000111) ? 48'b100100110111101101100010000100110111101101100010 :
(key == 11'b11011001000) ? 48'b100100110111000010000010000100110111000010000010 :
(key == 11'b11011001001) ? 48'b100100110110010110100101000100110110010110100101 :
(key == 11'b11011001010) ? 48'b100100110101101011001010000100110101101011001010 :
(key == 11'b11011001011) ? 48'b100100110100111111110010000100110100111111110010 :
(key == 11'b11011001100) ? 48'b100100110100010100011100000100110100010100011100 :
(key == 11'b11011001101) ? 48'b100100110011101001001001000100110011101001001001 :
(key == 11'b11011001110) ? 48'b100100110010111101111000000100110010111101111000 :
(key == 11'b11011001111) ? 48'b100100110010010010101010000100110010010010101010 :
(key == 11'b11011010000) ? 48'b100100110001100111011110000100110001100111011110 :
(key == 11'b11011010001) ? 48'b100100110000111100010100000100110000111100010100 :
(key == 11'b11011010010) ? 48'b100100110000010001001100000100110000010001001100 :
(key == 11'b11011010011) ? 48'b100100101111100110000110000100101111100110000110 :
(key == 11'b11011010100) ? 48'b100100101110111011000100000100101110111011000100 :
(key == 11'b11011010101) ? 48'b100100101110010000000100000100101110010000000100 :
(key == 11'b11011010110) ? 48'b100100101101100101000110000100101101100101000110 :
(key == 11'b11011010111) ? 48'b100100101100111010001010000100101100111010001010 :
(key == 11'b11011011000) ? 48'b100100101100001111010000000100101100001111010000 :
(key == 11'b11011011001) ? 48'b100100101011100100011010000100101011100100011010 :
(key == 11'b11011011010) ? 48'b100100101010111001100110000100101010111001100110 :
(key == 11'b11011011011) ? 48'b100100101010001110110010000100101010001110110010 :
(key == 11'b11011011100) ? 48'b100100101001100100000010000100101001100100000010 :
(key == 11'b11011011101) ? 48'b100100101000111001010110000100101000111001010110 :
(key == 11'b11011011110) ? 48'b100100101000001110101010000100101000001110101010 :
(key == 11'b11011011111) ? 48'b100100100111100100000000000100100111100100000000 :
(key == 11'b11011100000) ? 48'b100100100110111001011010000100100110111001011010 :
(key == 11'b11011100001) ? 48'b100100100110001110110101000100100110001110110101 :
(key == 11'b11011100010) ? 48'b100100100101100100010011000100100101100100010011 :
(key == 11'b11011100011) ? 48'b100100100100111001110100000100100100111001110100 :
(key == 11'b11011100100) ? 48'b100100100100001111010110000100100100001111010110 :
(key == 11'b11011100101) ? 48'b100100100011100100111100000100100011100100111100 :
(key == 11'b11011100110) ? 48'b100100100010111010100010000100100010111010100010 :
(key == 11'b11011100111) ? 48'b100100100010010000001100000100100010010000001100 :
(key == 11'b11011101000) ? 48'b100100100001100101111000000100100001100101111000 :
(key == 11'b11011101001) ? 48'b100100100000111011100110000100100000111011100110 :
(key == 11'b11011101010) ? 48'b100100100000010001010110000100100000010001010110 :
(key == 11'b11011101011) ? 48'b100100011111100111001001000100011111100111001001 :
(key == 11'b11011101100) ? 48'b100100011110111100111110000100011110111100111110 :
(key == 11'b11011101101) ? 48'b100100011110010010110101000100011110010010110101 :
(key == 11'b11011101110) ? 48'b100100011101101000101110000100011101101000101110 :
(key == 11'b11011101111) ? 48'b100100011100111110101011000100011100111110101011 :
(key == 11'b11011110000) ? 48'b100100011100010100101000000100011100010100101000 :
(key == 11'b11011110001) ? 48'b100100011011101010101001000100011011101010101001 :
(key == 11'b11011110010) ? 48'b100100011011000000101100000100011011000000101100 :
(key == 11'b11011110011) ? 48'b100100011010010110110010000100011010010110110010 :
(key == 11'b11011110100) ? 48'b100100011001101100111000000100011001101100111000 :
(key == 11'b11011110101) ? 48'b100100011001000011000001000100011001000011000001 :
(key == 11'b11011110110) ? 48'b100100011000011001001100000100011000011001001100 :
(key == 11'b11011110111) ? 48'b100100010111101111011100000100010111101111011100 :
(key == 11'b11011111000) ? 48'b100100010111000101101011000100010111000101101011 :
(key == 11'b11011111001) ? 48'b100100010110011011111101000100010110011011111101 :
(key == 11'b11011111010) ? 48'b100100010101110010010010000100010101110010010010 :
(key == 11'b11011111011) ? 48'b100100010101001000101010000100010101001000101010 :
(key == 11'b11011111100) ? 48'b100100010100011111000010000100010100011111000010 :
(key == 11'b11011111101) ? 48'b100100010011110101011101000100010011110101011101 :
(key == 11'b11011111110) ? 48'b100100010011001011111010000100010011001011111010 :
(key == 11'b11011111111) ? 48'b100100010010100010011100000100010010100010011100 :
(key == 11'b11100000000) ? 48'b100100010001111000111101000100010001111000111101 :
(key == 11'b11100000001) ? 48'b100100010001001111100001000100010001001111100001 :
(key == 11'b11100000010) ? 48'b100100010000100110001000000100010000100110001000 :
(key == 11'b11100000011) ? 48'b100100001111111100110000000100001111111100110000 :
(key == 11'b11100000100) ? 48'b100100001111010011011100000100001111010011011100 :
(key == 11'b11100000101) ? 48'b100100001110101010001000000100001110101010001000 :
(key == 11'b11100000110) ? 48'b100100001110000000111000000100001110000000111000 :
(key == 11'b11100000111) ? 48'b100100001101010111101001000100001101010111101001 :
(key == 11'b11100001000) ? 48'b100100001100101110011101000100001100101110011101 :
(key == 11'b11100001001) ? 48'b100100001100000101010011000100001100000101010011 :
(key == 11'b11100001010) ? 48'b100100001011011100001011000100001011011100001011 :
(key == 11'b11100001011) ? 48'b100100001010110011000101000100001010110011000101 :
(key == 11'b11100001100) ? 48'b100100001010001010000010000100001010001010000010 :
(key == 11'b11100001101) ? 48'b100100001001100001000000000100001001100001000000 :
(key == 11'b11100001110) ? 48'b100100001000111000000001000100001000111000000001 :
(key == 11'b11100001111) ? 48'b100100001000001111000100000100001000001111000100 :
(key == 11'b11100010000) ? 48'b100100000111100110001001000100000111100110001001 :
(key == 11'b11100010001) ? 48'b100100000110111101010001000100000110111101010001 :
(key == 11'b11100010010) ? 48'b100100000110010100011010000100000110010100011010 :
(key == 11'b11100010011) ? 48'b100100000101101011100110000100000101101011100110 :
(key == 11'b11100010100) ? 48'b100100000101000010110100000100000101000010110100 :
(key == 11'b11100010101) ? 48'b100100000100011010000100000100000100011010000100 :
(key == 11'b11100010110) ? 48'b100100000011110001010110000100000011110001010110 :
(key == 11'b11100010111) ? 48'b100100000011001000101010000100000011001000101010 :
(key == 11'b11100011000) ? 48'b100100000010100000000000000100000010100000000000 :
(key == 11'b11100011001) ? 48'b100100000001110111011001000100000001110111011001 :
(key == 11'b11100011010) ? 48'b100100000001001110110100000100000001001110110100 :
(key == 11'b11100011011) ? 48'b100100000000100110010010000100000000100110010010 :
(key == 11'b11100011100) ? 48'b100011111111111101110001000011111111111101110001 :
(key == 11'b11100011101) ? 48'b100011111111010101010010000011111111010101010010 :
(key == 11'b11100011110) ? 48'b100011111110101100110100000011111110101100110100 :
(key == 11'b11100011111) ? 48'b100011111110000100011010000011111110000100011010 :
(key == 11'b11100100000) ? 48'b100011111101011100000010000011111101011100000010 :
(key == 11'b11100100001) ? 48'b100011111100110011101011000011111100110011101011 :
(key == 11'b11100100010) ? 48'b100011111100001011010111000011111100001011010111 :
(key == 11'b11100100011) ? 48'b100011111011100011000101000011111011100011000101 :
(key == 11'b11100100100) ? 48'b100011111010111010110101000011111010111010110101 :
(key == 11'b11100100101) ? 48'b100011111010010010100111000011111010010010100111 :
(key == 11'b11100100110) ? 48'b100011111001101010011100000011111001101010011100 :
(key == 11'b11100100111) ? 48'b100011111001000010010010000011111001000010010010 :
(key == 11'b11100101000) ? 48'b100011111000011010001010000011111000011010001010 :
(key == 11'b11100101001) ? 48'b100011110111110010000110000011110111110010000110 :
(key == 11'b11100101010) ? 48'b100011110111001010000010000011110111001010000010 :
(key == 11'b11100101011) ? 48'b100011110110100010000001000011110110100010000001 :
(key == 11'b11100101100) ? 48'b100011110101111010000010000011110101111010000010 :
(key == 11'b11100101101) ? 48'b100011110101010010000101000011110101010010000101 :
(key == 11'b11100101110) ? 48'b100011110100101010001001000011110100101010001001 :
(key == 11'b11100101111) ? 48'b100011110100000010010001000011110100000010010001 :
(key == 11'b11100110000) ? 48'b100011110011011010011010000011110011011010011010 :
(key == 11'b11100110001) ? 48'b100011110010110010100110000011110010110010100110 :
(key == 11'b11100110010) ? 48'b100011110010001010110010000011110010001010110010 :
(key == 11'b11100110011) ? 48'b100011110001100011000010000011110001100011000010 :
(key == 11'b11100110100) ? 48'b100011110000111011010011000011110000111011010011 :
(key == 11'b11100110101) ? 48'b100011110000010011100111000011110000010011100111 :
(key == 11'b11100110110) ? 48'b100011101111101011111101000011101111101011111101 :
(key == 11'b11100110111) ? 48'b100011101111000100010100000011101111000100010100 :
(key == 11'b11100111000) ? 48'b100011101110011100101110000011101110011100101110 :
(key == 11'b11100111001) ? 48'b100011101101110101001010000011101101110101001010 :
(key == 11'b11100111010) ? 48'b100011101101001101101000000011101101001101101000 :
(key == 11'b11100111011) ? 48'b100011101100100110001000000011101100100110001000 :
(key == 11'b11100111100) ? 48'b100011101011111110101010000011101011111110101010 :
(key == 11'b11100111101) ? 48'b100011101011010111001110000011101011010111001110 :
(key == 11'b11100111110) ? 48'b100011101010101111110100000011101010101111110100 :
(key == 11'b11100111111) ? 48'b100011101010001000011100000011101010001000011100 :
(key == 11'b11101000000) ? 48'b100011101001100001000110000011101001100001000110 :
(key == 11'b11101000001) ? 48'b100011101000111001110011000011101000111001110011 :
(key == 11'b11101000010) ? 48'b100011101000010010100001000011101000010010100001 :
(key == 11'b11101000011) ? 48'b100011100111101011010000000011100111101011010000 :
(key == 11'b11101000100) ? 48'b100011100111000100000011000011100111000100000011 :
(key == 11'b11101000101) ? 48'b100011100110011100110111000011100110011100110111 :
(key == 11'b11101000110) ? 48'b100011100101110101101101000011100101110101101101 :
(key == 11'b11101000111) ? 48'b100011100101001110100110000011100101001110100110 :
(key == 11'b11101001000) ? 48'b100011100100100111100000000011100100100111100000 :
(key == 11'b11101001001) ? 48'b100011100100000000011100000011100100000000011100 :
(key == 11'b11101001010) ? 48'b100011100011011001011010000011100011011001011010 :
(key == 11'b11101001011) ? 48'b100011100010110010011010000011100010110010011010 :
(key == 11'b11101001100) ? 48'b100011100010001011011110000011100010001011011110 :
(key == 11'b11101001101) ? 48'b100011100001100100100010000011100001100100100010 :
(key == 11'b11101001110) ? 48'b100011100000111101101000000011100000111101101000 :
(key == 11'b11101001111) ? 48'b100011100000010110110000000011100000010110110000 :
(key == 11'b11101010000) ? 48'b100011011111101111111010000011011111101111111010 :
(key == 11'b11101010001) ? 48'b100011011111001001000111000011011111001001000111 :
(key == 11'b11101010010) ? 48'b100011011110100010010101000011011110100010010101 :
(key == 11'b11101010011) ? 48'b100011011101111011100110000011011101111011100110 :
(key == 11'b11101010100) ? 48'b100011011101010100111000000011011101010100111000 :
(key == 11'b11101010101) ? 48'b100011011100101110001100000011011100101110001100 :
(key == 11'b11101010110) ? 48'b100011011100000111100010000011011100000111100010 :
(key == 11'b11101010111) ? 48'b100011011011100000111010000011011011100000111010 :
(key == 11'b11101011000) ? 48'b100011011010111010010100000011011010111010010100 :
(key == 11'b11101011001) ? 48'b100011011010010011110001000011011010010011110001 :
(key == 11'b11101011010) ? 48'b100011011001101101001111000011011001101101001111 :
(key == 11'b11101011011) ? 48'b100011011001000110101111000011011001000110101111 :
(key == 11'b11101011100) ? 48'b100011011000100000010001000011011000100000010001 :
(key == 11'b11101011101) ? 48'b100011010111111001110101000011010111111001110101 :
(key == 11'b11101011110) ? 48'b100011010111010011011011000011010111010011011011 :
(key == 11'b11101011111) ? 48'b100011010110101101000011000011010110101101000011 :
(key == 11'b11101100000) ? 48'b100011010110000110101101000011010110000110101101 :
(key == 11'b11101100001) ? 48'b100011010101100000011001000011010101100000011001 :
(key == 11'b11101100010) ? 48'b100011010100111010000111000011010100111010000111 :
(key == 11'b11101100011) ? 48'b100011010100010011110110000011010100010011110110 :
(key == 11'b11101100100) ? 48'b100011010011101101101000000011010011101101101000 :
(key == 11'b11101100101) ? 48'b100011010011000111011100000011010011000111011100 :
(key == 11'b11101100110) ? 48'b100011010010100001010010000011010010100001010010 :
(key == 11'b11101100111) ? 48'b100011010001111011001001000011010001111011001001 :
(key == 11'b11101101000) ? 48'b100011010001010101000010000011010001010101000010 :
(key == 11'b11101101001) ? 48'b100011010000101110111110000011010000101110111110 :
(key == 11'b11101101010) ? 48'b100011010000001000111011000011010000001000111011 :
(key == 11'b11101101011) ? 48'b100011001111100010111001000011001111100010111001 :
(key == 11'b11101101100) ? 48'b100011001110111100111010000011001110111100111010 :
(key == 11'b11101101101) ? 48'b100011001110010110111110000011001110010110111110 :
(key == 11'b11101101110) ? 48'b100011001101110001000100000011001101110001000100 :
(key == 11'b11101101111) ? 48'b100011001101001011001010000011001101001011001010 :
(key == 11'b11101110000) ? 48'b100011001100100101010010000011001100100101010010 :
(key == 11'b11101110001) ? 48'b100011001011111111011101000011001011111111011101 :
(key == 11'b11101110010) ? 48'b100011001011011001101010000011001011011001101010 :
(key == 11'b11101110011) ? 48'b100011001010110011111000000011001010110011111000 :
(key == 11'b11101110100) ? 48'b100011001010001110001000000011001010001110001000 :
(key == 11'b11101110101) ? 48'b100011001001101000011010000011001001101000011010 :
(key == 11'b11101110110) ? 48'b100011001001000010101110000011001001000010101110 :
(key == 11'b11101110111) ? 48'b100011001000011101000100000011001000011101000100 :
(key == 11'b11101111000) ? 48'b100011000111110111011101000011000111110111011101 :
(key == 11'b11101111001) ? 48'b100011000111010001110110000011000111010001110110 :
(key == 11'b11101111010) ? 48'b100011000110101100010010000011000110101100010010 :
(key == 11'b11101111011) ? 48'b100011000110000110110000000011000110000110110000 :
(key == 11'b11101111100) ? 48'b100011000101100001010000000011000101100001010000 :
(key == 11'b11101111101) ? 48'b100011000100111011110001000011000100111011110001 :
(key == 11'b11101111110) ? 48'b100011000100010110010100000011000100010110010100 :
(key == 11'b11101111111) ? 48'b100011000011110000111000000011000011110000111000 :
(key == 11'b11110000000) ? 48'b100011000011001011100000000011000011001011100000 :
(key == 11'b11110000001) ? 48'b100011000010100110001000000011000010100110001000 :
(key == 11'b11110000010) ? 48'b100011000010000000110011000011000010000000110011 :
(key == 11'b11110000011) ? 48'b100011000001011011100000000011000001011011100000 :
(key == 11'b11110000100) ? 48'b100011000000110110001110000011000000110110001110 :
(key == 11'b11110000101) ? 48'b100011000000010000111111000011000000010000111111 :
(key == 11'b11110000110) ? 48'b100010111111101011110001000010111111101011110001 :
(key == 11'b11110000111) ? 48'b100010111111000110100100000010111111000110100100 :
(key == 11'b11110001000) ? 48'b100010111110100001011010000010111110100001011010 :
(key == 11'b11110001001) ? 48'b100010111101111100010010000010111101111100010010 :
(key == 11'b11110001010) ? 48'b100010111101010111001011000010111101010111001011 :
(key == 11'b11110001011) ? 48'b100010111100110010000111000010111100110010000111 :
(key == 11'b11110001100) ? 48'b100010111100001101000100000010111100001101000100 :
(key == 11'b11110001101) ? 48'b100010111011101000000100000010111011101000000100 :
(key == 11'b11110001110) ? 48'b100010111011000011000100000010111011000011000100 :
(key == 11'b11110001111) ? 48'b100010111010011110000111000010111010011110000111 :
(key == 11'b11110010000) ? 48'b100010111001111001001011000010111001111001001011 :
(key == 11'b11110010001) ? 48'b100010111001010100010010000010111001010100010010 :
(key == 11'b11110010010) ? 48'b100010111000101111011010000010111000101111011010 :
(key == 11'b11110010011) ? 48'b100010111000001010100100000010111000001010100100 :
(key == 11'b11110010100) ? 48'b100010110111100101110000000010110111100101110000 :
(key == 11'b11110010101) ? 48'b100010110111000000111110000010110111000000111110 :
(key == 11'b11110010110) ? 48'b100010110110011100001101000010110110011100001101 :
(key == 11'b11110010111) ? 48'b100010110101110111011110000010110101110111011110 :
(key == 11'b11110011000) ? 48'b100010110101010010110010000010110101010010110010 :
(key == 11'b11110011001) ? 48'b100010110100101110000110000010110100101110000110 :
(key == 11'b11110011010) ? 48'b100010110100001001011110000010110100001001011110 :
(key == 11'b11110011011) ? 48'b100010110011100100110110000010110011100100110110 :
(key == 11'b11110011100) ? 48'b100010110011000000010000000010110011000000010000 :
(key == 11'b11110011101) ? 48'b100010110010011011101101000010110010011011101101 :
(key == 11'b11110011110) ? 48'b100010110001110111001010000010110001110111001010 :
(key == 11'b11110011111) ? 48'b100010110001010010101011000010110001010010101011 :
(key == 11'b11110100000) ? 48'b100010110000101110001100000010110000101110001100 :
(key == 11'b11110100001) ? 48'b100010110000001001101111000010110000001001101111 :
(key == 11'b11110100010) ? 48'b100010101111100101010100000010101111100101010100 :
(key == 11'b11110100011) ? 48'b100010101111000000111011000010101111000000111011 :
(key == 11'b11110100100) ? 48'b100010101110011100100100000010101110011100100100 :
(key == 11'b11110100101) ? 48'b100010101101111000001110000010101101111000001110 :
(key == 11'b11110100110) ? 48'b100010101101010011111010000010101101010011111010 :
(key == 11'b11110100111) ? 48'b100010101100101111101000000010101100101111101000 :
(key == 11'b11110101000) ? 48'b100010101100001011011000000010101100001011011000 :
(key == 11'b11110101001) ? 48'b100010101011100111001010000010101011100111001010 :
(key == 11'b11110101010) ? 48'b100010101011000010111110000010101011000010111110 :
(key == 11'b11110101011) ? 48'b100010101010011110110100000010101010011110110100 :
(key == 11'b11110101100) ? 48'b100010101001111010101010000010101001111010101010 :
(key == 11'b11110101101) ? 48'b100010101001010110100011000010101001010110100011 :
(key == 11'b11110101110) ? 48'b100010101000110010011101000010101000110010011101 :
(key == 11'b11110101111) ? 48'b100010101000001110011001000010101000001110011001 :
(key == 11'b11110110000) ? 48'b100010100111101010010111000010100111101010010111 :
(key == 11'b11110110001) ? 48'b100010100111000110010111000010100111000110010111 :
(key == 11'b11110110010) ? 48'b100010100110100010011000000010100110100010011000 :
(key == 11'b11110110011) ? 48'b100010100101111110011100000010100101111110011100 :
(key == 11'b11110110100) ? 48'b100010100101011010100001000010100101011010100001 :
(key == 11'b11110110101) ? 48'b100010100100110110101000000010100100110110101000 :
(key == 11'b11110110110) ? 48'b100010100100010010110000000010100100010010110000 :
(key == 11'b11110110111) ? 48'b100010100011101110111010000010100011101110111010 :
(key == 11'b11110111000) ? 48'b100010100011001011000110000010100011001011000110 :
(key == 11'b11110111001) ? 48'b100010100010100111010100000010100010100111010100 :
(key == 11'b11110111010) ? 48'b100010100010000011100100000010100010000011100100 :
(key == 11'b11110111011) ? 48'b100010100001011111110100000010100001011111110100 :
(key == 11'b11110111100) ? 48'b100010100000111100001000000010100000111100001000 :
(key == 11'b11110111101) ? 48'b100010100000011000011100000010100000011000011100 :
(key == 11'b11110111110) ? 48'b100010011111110100110011000010011111110100110011 :
(key == 11'b11110111111) ? 48'b100010011111010001001011000010011111010001001011 :
(key == 11'b11111000000) ? 48'b100010011110101101100100000010011110101101100100 :
(key == 11'b11111000001) ? 48'b100010011110001010000000000010011110001010000000 :
(key == 11'b11111000010) ? 48'b100010011101100110011101000010011101100110011101 :
(key == 11'b11111000011) ? 48'b100010011101000010111100000010011101000010111100 :
(key == 11'b11111000100) ? 48'b100010011100011111011100000010011100011111011100 :
(key == 11'b11111000101) ? 48'b100010011011111011111111000010011011111011111111 :
(key == 11'b11111000110) ? 48'b100010011011011000100011000010011011011000100011 :
(key == 11'b11111000111) ? 48'b100010011010110101001000000010011010110101001000 :
(key == 11'b11111001000) ? 48'b100010011010010001110000000010011010010001110000 :
(key == 11'b11111001001) ? 48'b100010011001101110011010000010011001101110011010 :
(key == 11'b11111001010) ? 48'b100010011001001011000100000010011001001011000100 :
(key == 11'b11111001011) ? 48'b100010011000100111110000000010011000100111110000 :
(key == 11'b11111001100) ? 48'b100010011000000100011111000010011000000100011111 :
(key == 11'b11111001101) ? 48'b100010010111100001001111000010010111100001001111 :
(key == 11'b11111001110) ? 48'b100010010110111110000001000010010110111110000001 :
(key == 11'b11111001111) ? 48'b100010010110011010110101000010010110011010110101 :
(key == 11'b11111010000) ? 48'b100010010101110111101010000010010101110111101010 :
(key == 11'b11111010001) ? 48'b100010010101010100100001000010010101010100100001 :
(key == 11'b11111010010) ? 48'b100010010100110001011001000010010100110001011001 :
(key == 11'b11111010011) ? 48'b100010010100001110010011000010010100001110010011 :
(key == 11'b11111010100) ? 48'b100010010011101011001111000010010011101011001111 :
(key == 11'b11111010101) ? 48'b100010010011001000001100000010010011001000001100 :
(key == 11'b11111010110) ? 48'b100010010010100101001100000010010010100101001100 :
(key == 11'b11111010111) ? 48'b100010010010000010001100000010010010000010001100 :
(key == 11'b11111011000) ? 48'b100010010001011111010000000010010001011111010000 :
(key == 11'b11111011001) ? 48'b100010010000111100010100000010010000111100010100 :
(key == 11'b11111011010) ? 48'b100010010000011001011010000010010000011001011010 :
(key == 11'b11111011011) ? 48'b100010001111110110100001000010001111110110100001 :
(key == 11'b11111011100) ? 48'b100010001111010011101010000010001111010011101010 :
(key == 11'b11111011101) ? 48'b100010001110110000110100000010001110110000110100 :
(key == 11'b11111011110) ? 48'b100010001110001110000001000010001110001110000001 :
(key == 11'b11111011111) ? 48'b100010001101101011010000000010001101101011010000 :
(key == 11'b11111100000) ? 48'b100010001101001000100000000010001101001000100000 :
(key == 11'b11111100001) ? 48'b100010001100100101110001000010001100100101110001 :
(key == 11'b11111100010) ? 48'b100010001100000011000100000010001100000011000100 :
(key == 11'b11111100011) ? 48'b100010001011100000011001000010001011100000011001 :
(key == 11'b11111100100) ? 48'b100010001010111101110000000010001010111101110000 :
(key == 11'b11111100101) ? 48'b100010001010011011001000000010001010011011001000 :
(key == 11'b11111100110) ? 48'b100010001001111000100001000010001001111000100001 :
(key == 11'b11111100111) ? 48'b100010001001010101111100000010001001010101111100 :
(key == 11'b11111101000) ? 48'b100010001000110011011010000010001000110011011010 :
(key == 11'b11111101001) ? 48'b100010001000010000111000000010001000010000111000 :
(key == 11'b11111101010) ? 48'b100010000111101110011000000010000111101110011000 :
(key == 11'b11111101011) ? 48'b100010000111001011111010000010000111001011111010 :
(key == 11'b11111101100) ? 48'b100010000110101001011110000010000110101001011110 :
(key == 11'b11111101101) ? 48'b100010000110000111000011000010000110000111000011 :
(key == 11'b11111101110) ? 48'b100010000101100100101010000010000101100100101010 :
(key == 11'b11111101111) ? 48'b100010000101000010010011000010000101000010010011 :
(key == 11'b11111110000) ? 48'b100010000100011111111101000010000100011111111101 :
(key == 11'b11111110001) ? 48'b100010000011111101101000000010000011111101101000 :
(key == 11'b11111110010) ? 48'b100010000011011011010110000010000011011011010110 :
(key == 11'b11111110011) ? 48'b100010000010111001000100000010000010111001000100 :
(key == 11'b11111110100) ? 48'b100010000010010110110101000010000010010110110101 :
(key == 11'b11111110101) ? 48'b100010000001110100100111000010000001110100100111 :
(key == 11'b11111110110) ? 48'b100010000001010010011010000010000001010010011010 :
(key == 11'b11111110111) ? 48'b100010000000110000010000000010000000110000010000 :
(key == 11'b11111111000) ? 48'b100010000000001110001000000010000000001110001000 :
(key == 11'b11111111001) ? 48'b100001111111101100000000000001111111101100000000 :
(key == 11'b11111111010) ? 48'b100001111111001001111010000001111111001001111010 :
(key == 11'b11111111011) ? 48'b100001111110100111110110000001111110100111110110 :
(key == 11'b11111111100) ? 48'b100001111110000101110100000001111110000101110100 :
(key == 11'b11111111101) ? 48'b100001111101100011110010000001111101100011110010 :
(key == 11'b11111111110) ? 48'b100001111101000001110010000001111101000001110010 :
(key == 11'b11111111111) ? 48'b100001111100011111110101000001111100011111110101 : 48'd0;

endmodule

`default_nettype wire
