`default_nettype none

module finv
   ( input wire [31:0] x,
     output wire [31:0] y,
     output wire ovf);

   /* TODO: assumptions
    * - inputs and output are not unnormal numbers or NaN or +-inf 
    * - if e is 0, the number is interpreted as +0
    * - overflow and underflow are treated as the same for ovf wire
    * - when underflow, y will be 0
    */

   // split sequence to each subsequence
   wire xs;
   wire [7:0] xe;
   wire [22:0] xm;
   assign {xs, xe, xm} = x;

   // calc s
   wire s;
   assign s = xs;

   // calc e
   wire [7:0] e;
   assign e = (xm == 23'd0) ? 8'd254 - xe : 8'd253 - xe; 

   // calc m
   wire [22:0] m;
   wire [46:0] val;
   wire [10:0] key;
   wire [11:0] v;
   assign {key, v} = xm;
   // lookup table and get constant and grad
   finv_lookup_table lt(key, val);
   wire [24:0] constant;
   wire [24:0] grad;
   // constant supplements 1 at the MSB
   assign constant = {1'b1, val[46:24], 1'b0};
   assign grad = {1'b0, val[23:0]};
   wire [49:0] grad2; // length 49 = 25 + 25 - 1
   assign grad2 = {1'b1, xm, 1'b0} * grad;
   wire [24:0] tmp_m;
   assign tmp_m = constant - grad2[48:24];
   assign m = (xm == 23'd0) ? 23'd0 : tmp_m[22:0];

   assign y = {s, e, m};
   assign ovf = 0;

endmodule

module finv_lookup_table
   ( input wire [10:0] key,
     output wire [46:0] value);

   assign value =
(key == 11'b00000000000) ? 47'b11111111111000000000001111111111110000000000011 :
(key == 11'b00000000001) ? 47'b11111111101000000001001111111111010000000011011 :
(key == 11'b00000000010) ? 47'b11111111011000000011001111111110110000001001011 :
(key == 11'b00000000011) ? 47'b11111111001000000110001111111110010000010010011 :
(key == 11'b00000000100) ? 47'b11111110111000001010001111111101110000011110011 :
(key == 11'b00000000101) ? 47'b11111110101000001111001111111101010000101101010 :
(key == 11'b00000000110) ? 47'b11111110011000010101000111111100110000111111000 :
(key == 11'b00000000111) ? 47'b11111110001000011100000111111100010001010011111 :
(key == 11'b00000001000) ? 47'b11111101111000100100000111111011110001101011111 :
(key == 11'b00000001001) ? 47'b11111101101000101100111111111011010010000110100 :
(key == 11'b00000001010) ? 47'b11111101011000110110111111111010110010100100011 :
(key == 11'b00000001011) ? 47'b11111101001001000001110111111010010011000100111 :
(key == 11'b00000001100) ? 47'b11111100111001001101101111111001110011101000011 :
(key == 11'b00000001101) ? 47'b11111100101001011010100111111001010100001110111 :
(key == 11'b00000001110) ? 47'b11111100011001101000011111111000110100111000011 :
(key == 11'b00000001111) ? 47'b11111100001001110111010111111000010101100100111 :
(key == 11'b00000010000) ? 47'b11111011111010000111000111110111110110010100000 :
(key == 11'b00000010001) ? 47'b11111011101010010111111111110111010111000110010 :
(key == 11'b00000010010) ? 47'b11111011011010101001101111110110110111111011011 :
(key == 11'b00000010011) ? 47'b11111011001010111100011111110110011000110011010 :
(key == 11'b00000010100) ? 47'b11111010111011010000000111110101111001101110000 :
(key == 11'b00000010101) ? 47'b11111010101011100100110111110101011010101011111 :
(key == 11'b00000010110) ? 47'b11111010011011111010011111110100111011101100011 :
(key == 11'b00000010111) ? 47'b11111010001100010001000111110100011100101111111 :
(key == 11'b00000011000) ? 47'b11111001111100101000101111110011111101110110011 :
(key == 11'b00000011001) ? 47'b11111001101101000001001111110011011110111111011 :
(key == 11'b00000011010) ? 47'b11111001011101011010101111110011000000001011100 :
(key == 11'b00000011011) ? 47'b11111001001101110101001111110010100001011010011 :
(key == 11'b00000011100) ? 47'b11111000111110010000100111110010000010101100000 :
(key == 11'b00000011101) ? 47'b11111000101110101101000111110001100100000000111 :
(key == 11'b00000011110) ? 47'b11111000011111001010010111110001000101011000001 :
(key == 11'b00000011111) ? 47'b11111000001111101000101111110000100110110010100 :
(key == 11'b00000100000) ? 47'b11111000000000000111111111110000001000001111100 :
(key == 11'b00000100001) ? 47'b11110111110000101000001111101111101001101111100 :
(key == 11'b00000100010) ? 47'b11110111100001001001010111101111001011010010001 :
(key == 11'b00000100011) ? 47'b11110111010001101011011111101110101100110111101 :
(key == 11'b00000100100) ? 47'b11110111000010001110100111101110001110100000000 :
(key == 11'b00000100101) ? 47'b11110110110010110010100111101101110000001011001 :
(key == 11'b00000100110) ? 47'b11110110100011010111100111101101010001111001000 :
(key == 11'b00000100111) ? 47'b11110110010011111101011111101100110011101001101 :
(key == 11'b00000101000) ? 47'b11110110000100100100010111101100010101011101001 :
(key == 11'b00000101001) ? 47'b11110101110101001100000111101011110111010011010 :
(key == 11'b00000101010) ? 47'b11110101100101110100110111101011011001001100010 :
(key == 11'b00000101011) ? 47'b11110101010110011110100111101010111011001000001 :
(key == 11'b00000101100) ? 47'b11110101000111001001001111101010011101000110110 :
(key == 11'b00000101101) ? 47'b11110100110111110100101111101001111111000111111 :
(key == 11'b00000101110) ? 47'b11110100101000100001001111101001100001001011111 :
(key == 11'b00000101111) ? 47'b11110100011001001110100111101001000011010010101 :
(key == 11'b00000110000) ? 47'b11110100001001111100111111101000100101011100001 :
(key == 11'b00000110001) ? 47'b11110011111010101100010111101000000111101000100 :
(key == 11'b00000110010) ? 47'b11110011101011011100100111100111101001110111100 :
(key == 11'b00000110011) ? 47'b11110011011100001101101111100111001100001001001 :
(key == 11'b00000110100) ? 47'b11110011001100111111101111100110101110011101011 :
(key == 11'b00000110101) ? 47'b11110010111101110010110111100110010000110100101 :
(key == 11'b00000110110) ? 47'b11110010101110100110101111100101110011001110011 :
(key == 11'b00000110111) ? 47'b11110010011111011011100111100101010101101010111 :
(key == 11'b00000111000) ? 47'b11110010010000010001010111100100111000001010001 :
(key == 11'b00000111001) ? 47'b11110010000001001000000111100100011010101100001 :
(key == 11'b00000111010) ? 47'b11110001110001111111101111100011111101010000101 :
(key == 11'b00000111011) ? 47'b11110001100010111000001111100011011111110111111 :
(key == 11'b00000111100) ? 47'b11110001010011110001101111100011000010100001111 :
(key == 11'b00000111101) ? 47'b11110001000100101100000111100010100101001110100 :
(key == 11'b00000111110) ? 47'b11110000110101100111010111100010000111111101101 :
(key == 11'b00000111111) ? 47'b11110000100110100011100111100001101010101111101 :
(key == 11'b00001000000) ? 47'b11110000010111100000101111100001001101100100010 :
(key == 11'b00001000001) ? 47'b11110000001000011110101111100000110000011011100 :
(key == 11'b00001000010) ? 47'b11101111111001011101101111100000010011010101100 :
(key == 11'b00001000011) ? 47'b11101111101010011101011111011111110110010001111 :
(key == 11'b00001000100) ? 47'b11101111011011011110010111011111011001010001010 :
(key == 11'b00001000101) ? 47'b11101111001100011111111111011110111100010011000 :
(key == 11'b00001000110) ? 47'b11101110111101100010011111011110011111010111010 :
(key == 11'b00001000111) ? 47'b11101110101110100101111111011110000010011110011 :
(key == 11'b00001001000) ? 47'b11101110011111101010010111011101100101101000000 :
(key == 11'b00001001001) ? 47'b11101110010000101111100111011101001000110100010 :
(key == 11'b00001001010) ? 47'b11101110000001110101110111011100101100000011010 :
(key == 11'b00001001011) ? 47'b11101101110010111100110111011100001111010100100 :
(key == 11'b00001001100) ? 47'b11101101100100000100110111011011110010101000110 :
(key == 11'b00001001101) ? 47'b11101101010101001101101111011011010101111111011 :
(key == 11'b00001001110) ? 47'b11101101000110010111011111011010111001011000101 :
(key == 11'b00001001111) ? 47'b11101100110111100010000111011010011100110100011 :
(key == 11'b00001010000) ? 47'b11101100101000101101101111011010000000010010111 :
(key == 11'b00001010001) ? 47'b11101100011001111010000111011001100011110011110 :
(key == 11'b00001010010) ? 47'b11101100001011000111011111011001000111010111011 :
(key == 11'b00001010011) ? 47'b11101011111100010101100111011000101010111101011 :
(key == 11'b00001010100) ? 47'b11101011101101100100101111011000001110100110000 :
(key == 11'b00001010101) ? 47'b11101011011110110100101111010111110010010001010 :
(key == 11'b00001010110) ? 47'b11101011010000000101100111010111010101111111000 :
(key == 11'b00001010111) ? 47'b11101011000001010111010111010110111001101111011 :
(key == 11'b00001011000) ? 47'b11101010110010101001111111010110011101100010001 :
(key == 11'b00001011001) ? 47'b11101010100011111101011111010110000001010111100 :
(key == 11'b00001011010) ? 47'b11101010010101010001111111010101100101001111101 :
(key == 11'b00001011011) ? 47'b11101010000110100111001111010101001001001010000 :
(key == 11'b00001011100) ? 47'b11101001110111111101010111010100101101000110111 :
(key == 11'b00001011101) ? 47'b11101001101001010100010111010100010001000110010 :
(key == 11'b00001011110) ? 47'b11101001011010101100001111010011110101001000001 :
(key == 11'b00001011111) ? 47'b11101001001100000101000111010011011001001100111 :
(key == 11'b00001100000) ? 47'b11101000111101011110101111010010111101010011110 :
(key == 11'b00001100001) ? 47'b11101000101110111001001111010010100001011101010 :
(key == 11'b00001100010) ? 47'b11101000100000010100100111010010000101101001001 :
(key == 11'b00001100011) ? 47'b11101000010001110000110111010001101001110111100 :
(key == 11'b00001100100) ? 47'b11101000000011001101111111010001001110001000100 :
(key == 11'b00001100101) ? 47'b11100111110100101011111111010000110010011011111 :
(key == 11'b00001100110) ? 47'b11100111100110001010110111010000010110110001110 :
(key == 11'b00001100111) ? 47'b11100111010111101010100111001111111011001010010 :
(key == 11'b00001101000) ? 47'b11100111001001001011000111001111011111100100111 :
(key == 11'b00001101001) ? 47'b11100110111010101100100111001111000100000010010 :
(key == 11'b00001101010) ? 47'b11100110101100001110110111001110101000100001111 :
(key == 11'b00001101011) ? 47'b11100110011101110010000111001110001101000100001 :
(key == 11'b00001101100) ? 47'b11100110001111010110000111001101110001101000110 :
(key == 11'b00001101101) ? 47'b11100110000000111010111111001101010110001111110 :
(key == 11'b00001101110) ? 47'b11100101110010100000101111001100111010111001010 :
(key == 11'b00001101111) ? 47'b11100101100100000111001111001100011111100101000 :
(key == 11'b00001110000) ? 47'b11100101010101101110101111001100000100010011100 :
(key == 11'b00001110001) ? 47'b11100101000111010110111111001011101001000100010 :
(key == 11'b00001110010) ? 47'b11100100111001000000000111001011001101110111011 :
(key == 11'b00001110011) ? 47'b11100100101010101010000111001010110010101101000 :
(key == 11'b00001110100) ? 47'b11100100011100010100111111001010010111100101000 :
(key == 11'b00001110101) ? 47'b11100100001110000000100111001001111100011111011 :
(key == 11'b00001110110) ? 47'b11100011111111101101001111001001100001011100011 :
(key == 11'b00001110111) ? 47'b11100011110001011010100111001001000110011011100 :
(key == 11'b00001111000) ? 47'b11100011100011001000110111001000101011011101001 :
(key == 11'b00001111001) ? 47'b11100011010100110111110111001000010000100001000 :
(key == 11'b00001111010) ? 47'b11100011000110100111101111000111110101100111011 :
(key == 11'b00001111011) ? 47'b11100010111000011000011111000111011010110000001 :
(key == 11'b00001111100) ? 47'b11100010101010001010000111000110111111111011010 :
(key == 11'b00001111101) ? 47'b11100010011011111100011111000110100101001000110 :
(key == 11'b00001111110) ? 47'b11100010001101101111101111000110001010011000100 :
(key == 11'b00001111111) ? 47'b11100001111111100011110111000101101111101010110 :
(key == 11'b00010000000) ? 47'b11100001110001011000101111000101010100111111010 :
(key == 11'b00010000001) ? 47'b11100001100011001110100111000100111010010110011 :
(key == 11'b00010000010) ? 47'b11100001010101000101000111000100011111101111100 :
(key == 11'b00010000011) ? 47'b11100001000110111100100111000100000101001011010 :
(key == 11'b00010000100) ? 47'b11100000111000110100110111000011101010101001010 :
(key == 11'b00010000101) ? 47'b11100000101010101101110111000011010000001001011 :
(key == 11'b00010000110) ? 47'b11100000011100100111110111000010110101101100001 :
(key == 11'b00010000111) ? 47'b11100000001110100010100111000010011011010001001 :
(key == 11'b00010001000) ? 47'b11100000000000011110000111000010000000111000010 :
(key == 11'b00010001001) ? 47'b11011111110010011010011111000001100110100001111 :
(key == 11'b00010001010) ? 47'b11011111100100010111101111000001001100001101110 :
(key == 11'b00010001011) ? 47'b11011111010110010101101111000000110001111011111 :
(key == 11'b00010001100) ? 47'b11011111001000010100100111000000010111101100100 :
(key == 11'b00010001101) ? 47'b11011110111010010100001110111111111101011111010 :
(key == 11'b00010001110) ? 47'b11011110101100010100101110111111100011010100011 :
(key == 11'b00010001111) ? 47'b11011110011110010101111110111111001001001011101 :
(key == 11'b00010010000) ? 47'b11011110010000011000000110111110101111000101011 :
(key == 11'b00010010001) ? 47'b11011110000010011011000110111110010101000001011 :
(key == 11'b00010010010) ? 47'b11011101110100011110110110111101111010111111101 :
(key == 11'b00010010011) ? 47'b11011101100110100011010110111101100001000000001 :
(key == 11'b00010010100) ? 47'b11011101011000101000101110111101000111000010111 :
(key == 11'b00010010101) ? 47'b11011101001010101110111110111100101101001000001 :
(key == 11'b00010010110) ? 47'b11011100111100110101111110111100010011001111011 :
(key == 11'b00010010111) ? 47'b11011100101110111101101110111011111001011000111 :
(key == 11'b00010011000) ? 47'b11011100100001000110010110111011011111100100110 :
(key == 11'b00010011001) ? 47'b11011100010011001111101110111011000101110010110 :
(key == 11'b00010011010) ? 47'b11011100000101011001111110111010101100000011001 :
(key == 11'b00010011011) ? 47'b11011011110111100100111110111010010010010101110 :
(key == 11'b00010011100) ? 47'b11011011101001110000110110111001111000101010101 :
(key == 11'b00010011101) ? 47'b11011011011011111101011110111001011111000001101 :
(key == 11'b00010011110) ? 47'b11011011001110001010111110111001000101011011001 :
(key == 11'b00010011111) ? 47'b11011011000000011001000110111000101011110110011 :
(key == 11'b00010100000) ? 47'b11011010110010101000001110111000010010010100010 :
(key == 11'b00010100001) ? 47'b11011010100100110111111110110111111000110100001 :
(key == 11'b00010100010) ? 47'b11011010010111001000100110110111011111010110010 :
(key == 11'b00010100011) ? 47'b11011010001001011010000110110111000101111010111 :
(key == 11'b00010100100) ? 47'b11011001111011101100001110110110101100100001010 :
(key == 11'b00010100101) ? 47'b11011001101101111111001110110110010011001010000 :
(key == 11'b00010100110) ? 47'b11011001100000010011000110110101111001110101001 :
(key == 11'b00010100111) ? 47'b11011001010010100111100110110101100000100010001 :
(key == 11'b00010101000) ? 47'b11011001000100111100111110110101000111010001100 :
(key == 11'b00010101001) ? 47'b11011000110111010011001110110100101110000011010 :
(key == 11'b00010101010) ? 47'b11011000101001101010000110110100010100110110111 :
(key == 11'b00010101011) ? 47'b11011000011100000001110110110011111011101100110 :
(key == 11'b00010101100) ? 47'b11011000001110011010011110110011100010100101000 :
(key == 11'b00010101101) ? 47'b11011000000000110011101110110011001001011111001 :
(key == 11'b00010101110) ? 47'b11010111110011001101110110110010110000011011101 :
(key == 11'b00010101111) ? 47'b11010111100101101000101110110010010111011010010 :
(key == 11'b00010110000) ? 47'b11010111011000000100010110110001111110011011000 :
(key == 11'b00010110001) ? 47'b11010111001010100000110110110001100101011110000 :
(key == 11'b00010110010) ? 47'b11010110111100111101111110110001001100100010111 :
(key == 11'b00010110011) ? 47'b11010110101111011011111110110000110011101010001 :
(key == 11'b00010110100) ? 47'b11010110100001111010101110110000011010110011011 :
(key == 11'b00010110101) ? 47'b11010110010100011010010110110000000001111111000 :
(key == 11'b00010110110) ? 47'b11010110000110111010101110101111101001001100110 :
(key == 11'b00010110111) ? 47'b11010101111001011011101110101111010000011100010 :
(key == 11'b00010111000) ? 47'b11010101101011111101100110101110110111101110010 :
(key == 11'b00010111001) ? 47'b11010101011110100000001110101110011111000010001 :
(key == 11'b00010111010) ? 47'b11010101010001000011101110101110000110011000100 :
(key == 11'b00010111011) ? 47'b11010101000011100111110110101101101101110000101 :
(key == 11'b00010111100) ? 47'b11010100110110001100110110101101010101001011000 :
(key == 11'b00010111101) ? 47'b11010100101000110010100110101100111100100111101 :
(key == 11'b00010111110) ? 47'b11010100011011011001000110101100100100000110001 :
(key == 11'b00010111111) ? 47'b11010100001110000000010110101100001011100110111 :
(key == 11'b00011000000) ? 47'b11010100000000101000010110101011110011001001101 :
(key == 11'b00011000001) ? 47'b11010011110011010001000110101011011010101110011 :
(key == 11'b00011000010) ? 47'b11010011100101111010100110101011000010010101010 :
(key == 11'b00011000011) ? 47'b11010011011000100100111110101010101001111110100 :
(key == 11'b00011000100) ? 47'b11010011001011001111111110101010010001101001100 :
(key == 11'b00011000101) ? 47'b11010010111101111011110110101001111001010110110 :
(key == 11'b00011000110) ? 47'b11010010110000101000011110101001100001000110001 :
(key == 11'b00011000111) ? 47'b11010010100011010101101110101001001000110111010 :
(key == 11'b00011001000) ? 47'b11010010010110000011110110101000110000101010110 :
(key == 11'b00011001001) ? 47'b11010010001000110010101110101000011000100000010 :
(key == 11'b00011001010) ? 47'b11010001111011100010010110101000000000010111111 :
(key == 11'b00011001011) ? 47'b11010001101110010010101110100111101000010001100 :
(key == 11'b00011001100) ? 47'b11010001100001000011110110100111010000001101010 :
(key == 11'b00011001101) ? 47'b11010001010011110101101110100110111000001010111 :
(key == 11'b00011001110) ? 47'b11010001000110101000010110100110100000001010110 :
(key == 11'b00011001111) ? 47'b11010000111001011011101110100110001000001100100 :
(key == 11'b00011010000) ? 47'b11010000101100001111110110100101110000010000011 :
(key == 11'b00011010001) ? 47'b11010000011111000100101110100101011000010110010 :
(key == 11'b00011010010) ? 47'b11010000010001111010010110100101000000011110010 :
(key == 11'b00011010011) ? 47'b11010000000100110000100110100100101000101000000 :
(key == 11'b00011010100) ? 47'b11001111110111100111101110100100010000110100000 :
(key == 11'b00011010101) ? 47'b11001111101010011111100110100011111001000010000 :
(key == 11'b00011010110) ? 47'b11001111011101011000001110100011100001010010001 :
(key == 11'b00011010111) ? 47'b11001111010000010001011110100011001001100100000 :
(key == 11'b00011011000) ? 47'b11001111000011001011100110100010110001111000001 :
(key == 11'b00011011001) ? 47'b11001110110110000110010110100010011010001110000 :
(key == 11'b00011011010) ? 47'b11001110101001000001111110100010000010100110001 :
(key == 11'b00011011011) ? 47'b11001110011011111110001110100001101011000000001 :
(key == 11'b00011011100) ? 47'b11001110001110111011001110100001010011011100001 :
(key == 11'b00011011101) ? 47'b11001110000001111000111110100000111011111010001 :
(key == 11'b00011011110) ? 47'b11001101110100110111011110100000100100011010001 :
(key == 11'b00011011111) ? 47'b11001101100111110110101110100000001100111100010 :
(key == 11'b00011100000) ? 47'b11001101011010110110101110011111110101100000010 :
(key == 11'b00011100001) ? 47'b11001101001101110111010110011111011110000110001 :
(key == 11'b00011100010) ? 47'b11001101000000111000110110011111000110101110010 :
(key == 11'b00011100011) ? 47'b11001100110011111010111110011110101111011000000 :
(key == 11'b00011100100) ? 47'b11001100100110111101110110011110011000000011111 :
(key == 11'b00011100101) ? 47'b11001100011010000001011110011110000000110001110 :
(key == 11'b00011100110) ? 47'b11001100001101000101110110011101101001100001101 :
(key == 11'b00011100111) ? 47'b11001100000000001010110110011101010010010011011 :
(key == 11'b00011101000) ? 47'b11001011110011010000101110011100111011000111010 :
(key == 11'b00011101001) ? 47'b11001011100110010111001110011100100011111100111 :
(key == 11'b00011101010) ? 47'b11001011011001011110011110011100001100110100100 :
(key == 11'b00011101011) ? 47'b11001011001100100110010110011011110101101101111 :
(key == 11'b00011101100) ? 47'b11001010111111101111000110011011011110101001100 :
(key == 11'b00011101101) ? 47'b11001010110010111000011110011011000111100110111 :
(key == 11'b00011101110) ? 47'b11001010100110000010100110011010110000100110010 :
(key == 11'b00011101111) ? 47'b11001010011001001101011110011010011001100111101 :
(key == 11'b00011110000) ? 47'b11001010001100011000111110011010000010101010110 :
(key == 11'b00011110001) ? 47'b11001001111111100101001110011001101011101111111 :
(key == 11'b00011110010) ? 47'b11001001110010110010001110011001010100110111000 :
(key == 11'b00011110011) ? 47'b11001001100101111111111110011000111110000000001 :
(key == 11'b00011110100) ? 47'b11001001011001001110010110011000100111001010111 :
(key == 11'b00011110101) ? 47'b11001001001100011101011110011000010000010111110 :
(key == 11'b00011110110) ? 47'b11001000111111101101010110010111111001100110100 :
(key == 11'b00011110111) ? 47'b11001000110010111101110110010111100010110111001 :
(key == 11'b00011111000) ? 47'b11001000100110001111001110010111001100001001110 :
(key == 11'b00011111001) ? 47'b11001000011001100001000110010110110101011110000 :
(key == 11'b00011111010) ? 47'b11001000001100110011110110010110011110110100100 :
(key == 11'b00011111011) ? 47'b11001000000000000111001110010110001000001100110 :
(key == 11'b00011111100) ? 47'b11000111110011011011010110010101110001100110111 :
(key == 11'b00011111101) ? 47'b11000111100110110000000110010101011011000010110 :
(key == 11'b00011111110) ? 47'b11000111011010000101100110010101000100100000101 :
(key == 11'b00011111111) ? 47'b11000111001101011011110110010100101110000000011 :
(key == 11'b00100000000) ? 47'b11000111000000110010101110010100010111100010000 :
(key == 11'b00100000001) ? 47'b11000110110100001010010110010100000001000101100 :
(key == 11'b00100000010) ? 47'b11000110100111100010101110010011101010101011000 :
(key == 11'b00100000011) ? 47'b11000110011010111011101110010011010100010010001 :
(key == 11'b00100000100) ? 47'b11000110001110010101011110010010111101111011010 :
(key == 11'b00100000101) ? 47'b11000110000001101111110110010010100111100110010 :
(key == 11'b00100000110) ? 47'b11000101110101001010111110010010010001010011000 :
(key == 11'b00100000111) ? 47'b11000101101000100110101110010001111011000001101 :
(key == 11'b00100001000) ? 47'b11000101011100000011001110010001100100110010001 :
(key == 11'b00100001001) ? 47'b11000101001111100000011110010001001110100100100 :
(key == 11'b00100001010) ? 47'b11000101000010111110010110010000111000011000101 :
(key == 11'b00100001011) ? 47'b11000100110110011100111110010000100010001110110 :
(key == 11'b00100001100) ? 47'b11000100101001111100001110010000001100000110101 :
(key == 11'b00100001101) ? 47'b11000100011101011100001110001111110110000000011 :
(key == 11'b00100001110) ? 47'b11000100010000111100110110001111011111111011111 :
(key == 11'b00100001111) ? 47'b11000100000100011110001110001111001001111001010 :
(key == 11'b00100010000) ? 47'b11000011111000000000001110001110110011111000011 :
(key == 11'b00100010001) ? 47'b11000011101011100010111110001110011101111001011 :
(key == 11'b00100010010) ? 47'b11000011011111000110010110001110000111111100001 :
(key == 11'b00100010011) ? 47'b11000011010010101010011110001101110010000000111 :
(key == 11'b00100010100) ? 47'b11000011000110001111001110001101011100000111010 :
(key == 11'b00100010101) ? 47'b11000010111001110100101110001101000110001111100 :
(key == 11'b00100010110) ? 47'b11000010101101011010110110001100110000011001100 :
(key == 11'b00100010111) ? 47'b11000010100001000001100110001100011010100101010 :
(key == 11'b00100011000) ? 47'b11000010010100101001001110001100000100110011001 :
(key == 11'b00100011001) ? 47'b11000010001000010001010110001011101111000010100 :
(key == 11'b00100011010) ? 47'b11000001111011111010001110001011011001010011110 :
(key == 11'b00100011011) ? 47'b11000001101111100011101110001011000011100110101 :
(key == 11'b00100011100) ? 47'b11000001100011001101111110001010101101111011100 :
(key == 11'b00100011101) ? 47'b11000001010110111000110110001010011000010010000 :
(key == 11'b00100011110) ? 47'b11000001001010100100011110001010000010101010100 :
(key == 11'b00100011111) ? 47'b11000000111110010000101110001001101101000100101 :
(key == 11'b00100100000) ? 47'b11000000110001111101100110001001010111100000100 :
(key == 11'b00100100001) ? 47'b11000000100101101011001110001001000001111110010 :
(key == 11'b00100100010) ? 47'b11000000011001011001100110001000101100011101111 :
(key == 11'b00100100011) ? 47'b11000000001101001000011110001000010110111111000 :
(key == 11'b00100100100) ? 47'b11000000000000111000000110001000000001100010000 :
(key == 11'b00100100101) ? 47'b10111111110100101000010110000111101100000110110 :
(key == 11'b00100100110) ? 47'b10111111101000011001010110000111010110101101010 :
(key == 11'b00100100111) ? 47'b10111111011100001010111110000111000001010101100 :
(key == 11'b00100101000) ? 47'b10111111001111111101001110000110101011111111100 :
(key == 11'b00100101001) ? 47'b10111111000011110000001110000110010110101011010 :
(key == 11'b00100101010) ? 47'b10111110110111100011110110000110000001011000110 :
(key == 11'b00100101011) ? 47'b10111110101011011000000110000101101100001000000 :
(key == 11'b00100101100) ? 47'b10111110011111001101000110000101010110111001000 :
(key == 11'b00100101101) ? 47'b10111110010011000010101110000101000001101011110 :
(key == 11'b00100101110) ? 47'b10111110000110111000111110000100101100100000001 :
(key == 11'b00100101111) ? 47'b10111101111010101111111110000100010111010110100 :
(key == 11'b00100110000) ? 47'b10111101101110100111011110000100000010001110010 :
(key == 11'b00100110001) ? 47'b10111101100010011111101110000011101101000111110 :
(key == 11'b00100110010) ? 47'b10111101010110011000101110000011011000000011010 :
(key == 11'b00100110011) ? 47'b10111101001010010010001110000011000011000000010 :
(key == 11'b00100110100) ? 47'b10111100111110001100011110000010101101111111000 :
(key == 11'b00100110101) ? 47'b10111100110010000111010110000010011000111111100 :
(key == 11'b00100110110) ? 47'b10111100100110000010111110000010000100000001111 :
(key == 11'b00100110111) ? 47'b10111100011001111111000110000001101111000101101 :
(key == 11'b00100111000) ? 47'b10111100001101111011111110000001011010001011010 :
(key == 11'b00100111001) ? 47'b10111100000001111001011110000001000101010010100 :
(key == 11'b00100111010) ? 47'b10111011110101110111101110000000110000011011101 :
(key == 11'b00100111011) ? 47'b10111011101001110110011110000000011011100110010 :
(key == 11'b00100111100) ? 47'b10111011011101110101111110000000000110110010110 :
(key == 11'b00100111101) ? 47'b10111011010001110110000101111111110010000000111 :
(key == 11'b00100111110) ? 47'b10111011000101110110110101111111011101010000100 :
(key == 11'b00100111111) ? 47'b10111010111001111000001101111111001000100010000 :
(key == 11'b00101000000) ? 47'b10111010101101111010010101111110110011110101010 :
(key == 11'b00101000001) ? 47'b10111010100001111100111101111110011111001001111 :
(key == 11'b00101000010) ? 47'b10111010010110000000010101111110001010100000011 :
(key == 11'b00101000011) ? 47'b10111010001010000100010101111101110101111000100 :
(key == 11'b00101000100) ? 47'b10111001111110001000111101111101100001010010011 :
(key == 11'b00101000101) ? 47'b10111001110010001110001101111101001100101101110 :
(key == 11'b00101000110) ? 47'b10111001100110010100001101111100111000001011000 :
(key == 11'b00101000111) ? 47'b10111001011010011010101101111100100011101001110 :
(key == 11'b00101001000) ? 47'b10111001001110100001111101111100001111001010010 :
(key == 11'b00101001001) ? 47'b10111001000010101001110101111011111010101100011 :
(key == 11'b00101001010) ? 47'b10111000110110110010001101111011100110010000000 :
(key == 11'b00101001011) ? 47'b10111000101010111011010101111011010001110101011 :
(key == 11'b00101001100) ? 47'b10111000011111000101001101111010111101011100110 :
(key == 11'b00101001101) ? 47'b10111000010011001111100101111010101001000101011 :
(key == 11'b00101001110) ? 47'b10111000000111011010100101111010010100101111101 :
(key == 11'b00101001111) ? 47'b10110111111011100110001101111010000000011011101 :
(key == 11'b00101010000) ? 47'b10110111101111110010100101111001101100001001010 :
(key == 11'b00101010001) ? 47'b10110111100011111111011101111001010111111000100 :
(key == 11'b00101010010) ? 47'b10110111011000001101000101111001000011101001011 :
(key == 11'b00101010011) ? 47'b10110111001100011011001101111000101111011011111 :
(key == 11'b00101010100) ? 47'b10110111000000101010000101111000011011010000000 :
(key == 11'b00101010101) ? 47'b10110110110100111001100101111000000111000101111 :
(key == 11'b00101010110) ? 47'b10110110101001001001101101110111110010111101010 :
(key == 11'b00101010111) ? 47'b10110110011101011010010101110111011110110110001 :
(key == 11'b00101011000) ? 47'b10110110010001101011101101110111001010110000110 :
(key == 11'b00101011001) ? 47'b10110110000101111101101101110110110110101101000 :
(key == 11'b00101011010) ? 47'b10110101111010010000010101110110100010101010111 :
(key == 11'b00101011011) ? 47'b10110101101110100011100101110110001110101010011 :
(key == 11'b00101011100) ? 47'b10110101100010110111010101110101111010101011001 :
(key == 11'b00101011101) ? 47'b10110101010111001011110101110101100110101101111 :
(key == 11'b00101011110) ? 47'b10110101001011100000111101110101010010110010001 :
(key == 11'b00101011111) ? 47'b10110100111111110110101101110100111110111000000 :
(key == 11'b00101100000) ? 47'b10110100110100001101000101110100101010111111100 :
(key == 11'b00101100001) ? 47'b10110100101000100011111101110100010111001000011 :
(key == 11'b00101100010) ? 47'b10110100011100111011100101110100000011010011000 :
(key == 11'b00101100011) ? 47'b10110100010001010011110101110011101111011111010 :
(key == 11'b00101100100) ? 47'b10110100000101101100100101110011011011101100111 :
(key == 11'b00101100101) ? 47'b10110011111010000110000101110011000111111100010 :
(key == 11'b00101100110) ? 47'b10110011101110100000000101110010110100001101001 :
(key == 11'b00101100111) ? 47'b10110011100010111010110101110010100000011111110 :
(key == 11'b00101101000) ? 47'b10110011010111010110000101110010001100110011110 :
(key == 11'b00101101001) ? 47'b10110011001011110001111101110001111001001001010 :
(key == 11'b00101101010) ? 47'b10110011000000001110100101110001100101100000101 :
(key == 11'b00101101011) ? 47'b10110010110100101011101101110001010001111001011 :
(key == 11'b00101101100) ? 47'b10110010101001001001011101110000111110010011110 :
(key == 11'b00101101101) ? 47'b10110010011101100111101101110000101010101111011 :
(key == 11'b00101101110) ? 47'b10110010010010000110101101110000010111001100111 :
(key == 11'b00101101111) ? 47'b10110010000110100110010101110000000011101011111 :
(key == 11'b00101110000) ? 47'b10110001111011000110011101101111110000001100011 :
(key == 11'b00101110001) ? 47'b10110001101111100111010101101111011100101110101 :
(key == 11'b00101110010) ? 47'b10110001100100001000101101101111001001010010001 :
(key == 11'b00101110011) ? 47'b10110001011000101010101101101110110101110111010 :
(key == 11'b00101110100) ? 47'b10110001001101001101010101101110100010011110000 :
(key == 11'b00101110101) ? 47'b10110001000001110000100101101110001111000110010 :
(key == 11'b00101110110) ? 47'b10110000110110010100011101101101111011110000001 :
(key == 11'b00101110111) ? 47'b10110000101010111000110101101101101000011011011 :
(key == 11'b00101111000) ? 47'b10110000011111011101110101101101010101001000001 :
(key == 11'b00101111001) ? 47'b10110000010100000011011101101101000001110110100 :
(key == 11'b00101111010) ? 47'b10110000001000101001101101101100101110100110011 :
(key == 11'b00101111011) ? 47'b10101111111101010000100101101100011011010111111 :
(key == 11'b00101111100) ? 47'b10101111110001111000000101101100001000001010111 :
(key == 11'b00101111101) ? 47'b10101111100110100000000101101011110100111111010 :
(key == 11'b00101111110) ? 47'b10101111011011001000101101101011100001110101010 :
(key == 11'b00101111111) ? 47'b10101111001111110001111101101011001110101100110 :
(key == 11'b00110000000) ? 47'b10101111000100011011110101101010111011100101110 :
(key == 11'b00110000001) ? 47'b10101110111001000110001101101010101000100000001 :
(key == 11'b00110000010) ? 47'b10101110101101110001010101101010010101011100011 :
(key == 11'b00110000011) ? 47'b10101110100010011100111101101010000010011001111 :
(key == 11'b00110000100) ? 47'b10101110010111001001000101101001101111011000101 :
(key == 11'b00110000101) ? 47'b10101110001011110101111101101001011100011001010 :
(key == 11'b00110000110) ? 47'b10101110000000100011010101101001001001011011010 :
(key == 11'b00110000111) ? 47'b10101101110101010001010101101000110110011110110 :
(key == 11'b00110001000) ? 47'b10101101101001111111111101101000100011100011110 :
(key == 11'b00110001001) ? 47'b10101101011110101111000101101000010000101010001 :
(key == 11'b00110001010) ? 47'b10101101010011011110111101100111111101110010010 :
(key == 11'b00110001011) ? 47'b10101101001000001111010101100111101010111011110 :
(key == 11'b00110001100) ? 47'b10101100111101000000001101100111011000000110100 :
(key == 11'b00110001101) ? 47'b10101100110001110001101101100111000101010010110 :
(key == 11'b00110001110) ? 47'b10101100100110100011111101100110110010100000111 :
(key == 11'b00110001111) ? 47'b10101100011011010110100101100110011111110000001 :
(key == 11'b00110010000) ? 47'b10101100010000001001111101100110001101000001000 :
(key == 11'b00110010001) ? 47'b10101100000100111101110101100101111010010011010 :
(key == 11'b00110010010) ? 47'b10101011111001110010001101100101100111100110111 :
(key == 11'b00110010011) ? 47'b10101011101110100111010101100101010100111100010 :
(key == 11'b00110010100) ? 47'b10101011100011011100111101100101000010010010111 :
(key == 11'b00110010101) ? 47'b10101011011000010011001101100100101111101011000 :
(key == 11'b00110010110) ? 47'b10101011001101001001111101100100011101000100100 :
(key == 11'b00110010111) ? 47'b10101011000010000001010101100100001010011111101 :
(key == 11'b00110011000) ? 47'b10101010110110111001010101100011110111111100001 :
(key == 11'b00110011001) ? 47'b10101010101011110001110101100011100101011010000 :
(key == 11'b00110011010) ? 47'b10101010100000101010111101100011010010111001011 :
(key == 11'b00110011011) ? 47'b10101010010101100100101101100011000000011010011 :
(key == 11'b00110011100) ? 47'b10101010001010011110111101100010101101111100101 :
(key == 11'b00110011101) ? 47'b10101001111111011001110101100010011011100000011 :
(key == 11'b00110011110) ? 47'b10101001110100010101001101100010001001000101011 :
(key == 11'b00110011111) ? 47'b10101001101001010001001101100001110110101100000 :
(key == 11'b00110100000) ? 47'b10101001011110001101110101100001100100010100001 :
(key == 11'b00110100001) ? 47'b10101001010011001010111101100001010001111101100 :
(key == 11'b00110100010) ? 47'b10101001001000001000101101100000111111101000100 :
(key == 11'b00110100011) ? 47'b10101000111101000110111101100000101101010100101 :
(key == 11'b00110100100) ? 47'b10101000110010000101110101100000011011000010011 :
(key == 11'b00110100101) ? 47'b10101000100111000101010101100000001000110001101 :
(key == 11'b00110100110) ? 47'b10101000011100000101010101011111110110100010010 :
(key == 11'b00110100111) ? 47'b10101000010001000101111101011111100100010100010 :
(key == 11'b00110101000) ? 47'b10101000000110000111000101011111010010000111101 :
(key == 11'b00110101001) ? 47'b10100111111011001000101101011110111111111100011 :
(key == 11'b00110101010) ? 47'b10100111110000001011000101011110101101110010110 :
(key == 11'b00110101011) ? 47'b10100111100101001101111101011110011011101010011 :
(key == 11'b00110101100) ? 47'b10100111011010010001010101011110001001100011011 :
(key == 11'b00110101101) ? 47'b10100111001111010101010101011101110111011101111 :
(key == 11'b00110101110) ? 47'b10100111000100011001110101011101100101011001101 :
(key == 11'b00110101111) ? 47'b10100110111001011110111101011101010011010110111 :
(key == 11'b00110110000) ? 47'b10100110101110100100100101011101000001010101011 :
(key == 11'b00110110001) ? 47'b10100110100011101010110101011100101111010101100 :
(key == 11'b00110110010) ? 47'b10100110011000110001101101011100011101010111000 :
(key == 11'b00110110011) ? 47'b10100110001101111001000101011100001011011001111 :
(key == 11'b00110110100) ? 47'b10100110000011000000111101011011111001011110000 :
(key == 11'b00110110101) ? 47'b10100101111000001001011101011011100111100011101 :
(key == 11'b00110110110) ? 47'b10100101101101010010011101011011010101101010100 :
(key == 11'b00110110111) ? 47'b10100101100010011100000101011011000011110010111 :
(key == 11'b00110111000) ? 47'b10100101010111100110001101011010110001111100100 :
(key == 11'b00110111001) ? 47'b10100101001100110000111101011010100000000111110 :
(key == 11'b00110111010) ? 47'b10100101000001111100001101011010001110010100001 :
(key == 11'b00110111011) ? 47'b10100100110111001000000101011001111100100010000 :
(key == 11'b00110111100) ? 47'b10100100101100010100011101011001101010110001010 :
(key == 11'b00110111101) ? 47'b10100100100001100001011101011001011001000010000 :
(key == 11'b00110111110) ? 47'b10100100010110101110111101011001000111010011111 :
(key == 11'b00110111111) ? 47'b10100100001011111100111101011000110101100111001 :
(key == 11'b00111000000) ? 47'b10100100000001001011100101011000100011111011111 :
(key == 11'b00111000001) ? 47'b10100011110110011010101101011000010010010001111 :
(key == 11'b00111000010) ? 47'b10100011101011101010011101011000000000101001011 :
(key == 11'b00111000011) ? 47'b10100011100000111010101101010111101111000010001 :
(key == 11'b00111000100) ? 47'b10100011010110001011011101010111011101011100001 :
(key == 11'b00111000101) ? 47'b10100011001011011100110101010111001011110111100 :
(key == 11'b00111000110) ? 47'b10100011000000101110101101010110111010010100011 :
(key == 11'b00111000111) ? 47'b10100010110110000001001101010110101000110010100 :
(key == 11'b00111001000) ? 47'b10100010101011010100001101010110010111010010000 :
(key == 11'b00111001001) ? 47'b10100010100000100111101101010110000101110010110 :
(key == 11'b00111001010) ? 47'b10100010010101111011110101010101110100010101000 :
(key == 11'b00111001011) ? 47'b10100010001011010000011101010101100010111000100 :
(key == 11'b00111001100) ? 47'b10100010000000100101100101010101010001011101010 :
(key == 11'b00111001101) ? 47'b10100001110101111011010101010101000000000011100 :
(key == 11'b00111001110) ? 47'b10100001101011010001100101010100101110101010111 :
(key == 11'b00111001111) ? 47'b10100001100000101000011101010100011101010011111 :
(key == 11'b00111010000) ? 47'b10100001010101111111110101010100001011111110000 :
(key == 11'b00111010001) ? 47'b10100001001011010111101101010011111010101001100 :
(key == 11'b00111010010) ? 47'b10100001000000110000000101010011101001010110010 :
(key == 11'b00111010011) ? 47'b10100000110110001001000101010011011000000100011 :
(key == 11'b00111010100) ? 47'b10100000101011100010100101010011000110110011110 :
(key == 11'b00111010101) ? 47'b10100000100000111100101101010010110101100100101 :
(key == 11'b00111010110) ? 47'b10100000010110010111010101010010100100010110110 :
(key == 11'b00111010111) ? 47'b10100000001011110010011101010010010011001010001 :
(key == 11'b00111011000) ? 47'b10100000000001001110000101010010000001111110110 :
(key == 11'b00111011001) ? 47'b10011111110110101010010101010001110000110100111 :
(key == 11'b00111011010) ? 47'b10011111101100000111000101010001011111101100001 :
(key == 11'b00111011011) ? 47'b10011111100001100100010101010001001110100100110 :
(key == 11'b00111011100) ? 47'b10011111010111000010000101010000111101011110100 :
(key == 11'b00111011101) ? 47'b10011111001100100000011101010000101100011001110 :
(key == 11'b00111011110) ? 47'b10011111000001111111010101010000011011010110010 :
(key == 11'b00111011111) ? 47'b10011110110111011110101101010000001010010100000 :
(key == 11'b00111100000) ? 47'b10011110101100111110101101001111111001010011010 :
(key == 11'b00111100001) ? 47'b10011110100010011111001101001111101000010011101 :
(key == 11'b00111100010) ? 47'b10011110011000000000001101001111010111010101011 :
(key == 11'b00111100011) ? 47'b10011110001101100001101101001111000110011000010 :
(key == 11'b00111100100) ? 47'b10011110000011000011110101001110110101011100101 :
(key == 11'b00111100101) ? 47'b10011101111000100110010101001110100100100010000 :
(key == 11'b00111100110) ? 47'b10011101101110001001011101001110010011101000110 :
(key == 11'b00111100111) ? 47'b10011101100011101101001101001110000010110001000 :
(key == 11'b00111101000) ? 47'b10011101011001010001010101001101110001111010011 :
(key == 11'b00111101001) ? 47'b10011101001110110110000101001101100001000101000 :
(key == 11'b00111101010) ? 47'b10011101000100011011001101001101010000010000110 :
(key == 11'b00111101011) ? 47'b10011100111010000000111101001100111111011110000 :
(key == 11'b00111101100) ? 47'b10011100101111100111010101001100101110101100101 :
(key == 11'b00111101101) ? 47'b10011100100101001110000101001100011101111100010 :
(key == 11'b00111101110) ? 47'b10011100011010110101011101001100001101001101010 :
(key == 11'b00111101111) ? 47'b10011100010000011101010101001011111100011111101 :
(key == 11'b00111110000) ? 47'b10011100000110000101100101001011101011110010111 :
(key == 11'b00111110001) ? 47'b10011011111011101110100101001011011011000111111 :
(key == 11'b00111110010) ? 47'b10011011110001010111111101001011001010011101111 :
(key == 11'b00111110011) ? 47'b10011011100111000001110101001010111001110101000 :
(key == 11'b00111110100) ? 47'b10011011011100101100010101001010101001001101101 :
(key == 11'b00111110101) ? 47'b10011011010010010111010101001010011000100111100 :
(key == 11'b00111110110) ? 47'b10011011001000000010110101001010001000000010100 :
(key == 11'b00111110111) ? 47'b10011010111101101110110101001001110111011110111 :
(key == 11'b00111111000) ? 47'b10011010110011011011010101001001100110111100010 :
(key == 11'b00111111001) ? 47'b10011010101001001000010101001001010110011011000 :
(key == 11'b00111111010) ? 47'b10011010011110110101111101001001000101111011001 :
(key == 11'b00111111011) ? 47'b10011010010100100011111101001000110101011100010 :
(key == 11'b00111111100) ? 47'b10011010001010010010100101001000100100111110111 :
(key == 11'b00111111101) ? 47'b10011010000000000001101101001000010100100010101 :
(key == 11'b00111111110) ? 47'b10011001110101110001010101001000000100000111101 :
(key == 11'b00111111111) ? 47'b10011001101011100001011101000111110011101101110 :
(key == 11'b01000000000) ? 47'b10011001100001010010000101000111100011010101001 :
(key == 11'b01000000001) ? 47'b10011001010111000011001101000111010010111101110 :
(key == 11'b01000000010) ? 47'b10011001001100110100110101000111000010100111101 :
(key == 11'b01000000011) ? 47'b10011001000010100111000101000110110010010010111 :
(key == 11'b01000000100) ? 47'b10011000111000011001101101000110100001111111000 :
(key == 11'b01000000101) ? 47'b10011000101110001100111101000110010001101100110 :
(key == 11'b01000000110) ? 47'b10011000100100000000100101000110000001011011011 :
(key == 11'b01000000111) ? 47'b10011000011001110100110101000101110001001011011 :
(key == 11'b01000001000) ? 47'b10011000001111101001100101000101100000111100101 :
(key == 11'b01000001001) ? 47'b10011000000101011110110101000101010000101111001 :
(key == 11'b01000001010) ? 47'b10010111111011010100011101000101000000100010100 :
(key == 11'b01000001011) ? 47'b10010111110001001010101101000100110000010111011 :
(key == 11'b01000001100) ? 47'b10010111100111000001011101000100100000001101011 :
(key == 11'b01000001101) ? 47'b10010111011100111000101101000100010000000100101 :
(key == 11'b01000001110) ? 47'b10010111010010110000011101000011111111111101001 :
(key == 11'b01000001111) ? 47'b10010111001000101000101101000011101111110110110 :
(key == 11'b01000010000) ? 47'b10010110111110100001011101000011011111110001101 :
(key == 11'b01000010001) ? 47'b10010110110100011010101101000011001111101101101 :
(key == 11'b01000010010) ? 47'b10010110101010010100011101000010111111101010110 :
(key == 11'b01000010011) ? 47'b10010110100000001110110101000010101111101001011 :
(key == 11'b01000010100) ? 47'b10010110010110001001100101000010011111101001000 :
(key == 11'b01000010101) ? 47'b10010110001100000100110101000010001111101001111 :
(key == 11'b01000010110) ? 47'b10010110000010000000100101000001111111101011110 :
(key == 11'b01000010111) ? 47'b10010101110111111100110101000001101111101111000 :
(key == 11'b01000011000) ? 47'b10010101101101111001100101000001011111110011011 :
(key == 11'b01000011001) ? 47'b10010101100011110110110101000001001111111000111 :
(key == 11'b01000011010) ? 47'b10010101011001110100100101000000111111111111101 :
(key == 11'b01000011011) ? 47'b10010101001111110010110101000000110000000111100 :
(key == 11'b01000011100) ? 47'b10010101000101110001100101000000100000010000101 :
(key == 11'b01000011101) ? 47'b10010100111011110000110101000000010000011010111 :
(key == 11'b01000011110) ? 47'b10010100110001110000100101000000000000100110011 :
(key == 11'b01000011111) ? 47'b10010100100111110000110100111111110000110011000 :
(key == 11'b01000100000) ? 47'b10010100011101110001011100111111100001000000101 :
(key == 11'b01000100001) ? 47'b10010100010011110010101100111111010001001111101 :
(key == 11'b01000100010) ? 47'b10010100001001110100011100111111000001011111111 :
(key == 11'b01000100011) ? 47'b10010011111111110110100100111110110001110001000 :
(key == 11'b01000100100) ? 47'b10010011110101111001010100111110100010000011100 :
(key == 11'b01000100101) ? 47'b10010011101011111100011100111110010010010111001 :
(key == 11'b01000100110) ? 47'b10010011100010000000001100111110000010101100000 :
(key == 11'b01000100111) ? 47'b10010011011000000100010100111101110011000001111 :
(key == 11'b01000101000) ? 47'b10010011001110001000111100111101100011011000111 :
(key == 11'b01000101001) ? 47'b10010011000100001110000100111101010011110001001 :
(key == 11'b01000101010) ? 47'b10010010111010010011101100111101000100001010100 :
(key == 11'b01000101011) ? 47'b10010010110000011001110100111100110100100101000 :
(key == 11'b01000101100) ? 47'b10010010100110100000011100111100100101000000110 :
(key == 11'b01000101101) ? 47'b10010010011100100111100100111100010101011101101 :
(key == 11'b01000101110) ? 47'b10010010010010101111000100111100000101111011100 :
(key == 11'b01000101111) ? 47'b10010010001000110111001100111011110110011010110 :
(key == 11'b01000110000) ? 47'b10010001111110111111101100111011100110111010111 :
(key == 11'b01000110001) ? 47'b10010001110101001000101100111011010111011100010 :
(key == 11'b01000110010) ? 47'b10010001101011010010001100111011000111111110110 :
(key == 11'b01000110011) ? 47'b10010001100001011100001100111010111000100010100 :
(key == 11'b01000110100) ? 47'b10010001010111100110101100111010101001000111011 :
(key == 11'b01000110101) ? 47'b10010001001101110001101100111010011001101101011 :
(key == 11'b01000110110) ? 47'b10010001000011111101000100111010001010010100011 :
(key == 11'b01000110111) ? 47'b10010000111010001000111100111001111010111100100 :
(key == 11'b01000111000) ? 47'b10010000110000010101011100111001101011100110000 :
(key == 11'b01000111001) ? 47'b10010000100110100010010100111001011100010000011 :
(key == 11'b01000111010) ? 47'b10010000011100101111101100111001001100111100000 :
(key == 11'b01000111011) ? 47'b10010000010010111101011100111000111101101000101 :
(key == 11'b01000111100) ? 47'b10010000001001001011110100111000101110010110100 :
(key == 11'b01000111101) ? 47'b10001111111111011010100100111000011111000101011 :
(key == 11'b01000111110) ? 47'b10001111110101101001110100111000001111110101100 :
(key == 11'b01000111111) ? 47'b10001111101011111001100100111000000000100110101 :
(key == 11'b01001000000) ? 47'b10001111100010001001110100110111110001011001000 :
(key == 11'b01001000001) ? 47'b10001111011000011010011100110111100010001100010 :
(key == 11'b01001000010) ? 47'b10001111001110101011101100110111010011000000111 :
(key == 11'b01001000011) ? 47'b10001111000100111101010100110111000011110110100 :
(key == 11'b01001000100) ? 47'b10001110111011001111011100110110110100101101010 :
(key == 11'b01001000101) ? 47'b10001110110001100010000100110110100101100101001 :
(key == 11'b01001000110) ? 47'b10001110100111110101000100110110010110011110000 :
(key == 11'b01001000111) ? 47'b10001110011110001000100100110110000111011000000 :
(key == 11'b01001001000) ? 47'b10001110010100011100100100110101111000010011001 :
(key == 11'b01001001001) ? 47'b10001110001010110001000100110101101001001111011 :
(key == 11'b01001001010) ? 47'b10001110000001000110000100110101011010001100111 :
(key == 11'b01001001011) ? 47'b10001101110111011011011100110101001011001011010 :
(key == 11'b01001001100) ? 47'b10001101101101110001010100110100111100001010110 :
(key == 11'b01001001101) ? 47'b10001101100100000111101100110100101101001011011 :
(key == 11'b01001001110) ? 47'b10001101011010011110100100110100011110001101001 :
(key == 11'b01001001111) ? 47'b10001101010000110101110100110100001111001111111 :
(key == 11'b01001010000) ? 47'b10001101000111001101100100110100000000010011110 :
(key == 11'b01001010001) ? 47'b10001100111101100101110100110011110001011000110 :
(key == 11'b01001010010) ? 47'b10001100110011111110011100110011100010011110110 :
(key == 11'b01001010011) ? 47'b10001100101010010111100100110011010011100101111 :
(key == 11'b01001010100) ? 47'b10001100100000110001001100110011000100101110001 :
(key == 11'b01001010101) ? 47'b10001100010111001011010100110010110101110111100 :
(key == 11'b01001010110) ? 47'b10001100001101100101110100110010100111000001110 :
(key == 11'b01001010111) ? 47'b10001100000100000000111100110010011000001101011 :
(key == 11'b01001011000) ? 47'b10001011111010011100010100110010001001011001110 :
(key == 11'b01001011001) ? 47'b10001011110000111000010100110001111010100111100 :
(key == 11'b01001011010) ? 47'b10001011100111010100101100110001101011110110001 :
(key == 11'b01001011011) ? 47'b10001011011101110001100100110001011101000101111 :
(key == 11'b01001011100) ? 47'b10001011010100001110111100110001001110010110110 :
(key == 11'b01001011101) ? 47'b10001011001010101100101100110000111111101000101 :
(key == 11'b01001011110) ? 47'b10001011000001001010111100110000110000111011100 :
(key == 11'b01001011111) ? 47'b10001010110111101001100100110000100010001111011 :
(key == 11'b01001100000) ? 47'b10001010101110001000110100110000010011100100101 :
(key == 11'b01001100001) ? 47'b10001010100100101000011100110000000100111010110 :
(key == 11'b01001100010) ? 47'b10001010011011001000011100101111110110010001111 :
(key == 11'b01001100011) ? 47'b10001010010001101000111100101111100111101010000 :
(key == 11'b01001100100) ? 47'b10001010001000001001111100101111011001000011011 :
(key == 11'b01001100101) ? 47'b10001001111110101011011100101111001010011101110 :
(key == 11'b01001100110) ? 47'b10001001110101001101010100101110111011111001001 :
(key == 11'b01001100111) ? 47'b10001001101011101111101100101110101101010101101 :
(key == 11'b01001101000) ? 47'b10001001100010010010011100101110011110110011000 :
(key == 11'b01001101001) ? 47'b10001001011000110101101100101110010000010001100 :
(key == 11'b01001101010) ? 47'b10001001001111011001011100101110000001110001001 :
(key == 11'b01001101011) ? 47'b10001001000101111101101100101101110011010001111 :
(key == 11'b01001101100) ? 47'b10001000111100100010010100101101100100110011101 :
(key == 11'b01001101101) ? 47'b10001000110011000111010100101101010110010110010 :
(key == 11'b01001101110) ? 47'b10001000101001101100110100101101000111111001111 :
(key == 11'b01001101111) ? 47'b10001000100000010010110100101100111001011110110 :
(key == 11'b01001110000) ? 47'b10001000010110111001010100101100101011000100110 :
(key == 11'b01001110001) ? 47'b10001000001101100000001100101100011100101011100 :
(key == 11'b01001110010) ? 47'b10001000000100000111011100101100001110010011011 :
(key == 11'b01001110011) ? 47'b10000111111010101111010100101011111111111100011 :
(key == 11'b01001110100) ? 47'b10000111110001010111011100101011110001100110010 :
(key == 11'b01001110101) ? 47'b10000111101000000000001100101011100011010001011 :
(key == 11'b01001110110) ? 47'b10000111011110101001010100101011010100111101011 :
(key == 11'b01001110111) ? 47'b10000111010101010010110100101011000110101010010 :
(key == 11'b01001111000) ? 47'b10000111001011111100110100101010111000011000011 :
(key == 11'b01001111001) ? 47'b10000111000010100111010100101010101010000111100 :
(key == 11'b01001111010) ? 47'b10000110111001010010001100101010011011110111100 :
(key == 11'b01001111011) ? 47'b10000110101111111101100100101010001101101000101 :
(key == 11'b01001111100) ? 47'b10000110100110101001011100101001111111011011000 :
(key == 11'b01001111101) ? 47'b10000110011101010101100100101001110001001101111 :
(key == 11'b01001111110) ? 47'b10000110010100000010010100101001100011000010010 :
(key == 11'b01001111111) ? 47'b10000110001010101111011100101001010100110111011 :
(key == 11'b01010000000) ? 47'b10000110000001011100111100101001000110101101100 :
(key == 11'b01010000001) ? 47'b10000101111000001011000100101000111000100100111 :
(key == 11'b01010000010) ? 47'b10000101101110111001011100101000101010011101000 :
(key == 11'b01010000011) ? 47'b10000101100101101000010100101000011100010110001 :
(key == 11'b01010000100) ? 47'b10000101011100010111101100101000001110010000100 :
(key == 11'b01010000101) ? 47'b10000101010011000111011100101000000000001011101 :
(key == 11'b01010000110) ? 47'b10000101001001110111101100100111110010001000000 :
(key == 11'b01010000111) ? 47'b10000101000000101000010100100111100100000101001 :
(key == 11'b01010001000) ? 47'b10000100110111011001011100100111010110000011100 :
(key == 11'b01010001001) ? 47'b10000100101110001010111100100111001000000010101 :
(key == 11'b01010001010) ? 47'b10000100100100111100111100100110111010000010111 :
(key == 11'b01010001011) ? 47'b10000100011011101111010100100110101100000100001 :
(key == 11'b01010001100) ? 47'b10000100010010100010001100100110011110000110011 :
(key == 11'b01010001101) ? 47'b10000100001001010101011100100110010000001001101 :
(key == 11'b01010001110) ? 47'b10000100000000001001001100100110000010001101111 :
(key == 11'b01010001111) ? 47'b10000011110110111101010100100101110100010011000 :
(key == 11'b01010010000) ? 47'b10000011101101110001111100100101100110011001010 :
(key == 11'b01010010001) ? 47'b10000011100100100110111100100101011000100000011 :
(key == 11'b01010010010) ? 47'b10000011011011011100010100100101001010101000011 :
(key == 11'b01010010011) ? 47'b10000011010010010010001100100100111100110001100 :
(key == 11'b01010010100) ? 47'b10000011001001001000100100100100101110111011110 :
(key == 11'b01010010101) ? 47'b10000010111111111111010100100100100001000110111 :
(key == 11'b01010010110) ? 47'b10000010110110110110011100100100010011010010111 :
(key == 11'b01010010111) ? 47'b10000010101101101110000100100100000101100000000 :
(key == 11'b01010011000) ? 47'b10000010100100100110001100100011110111101110001 :
(key == 11'b01010011001) ? 47'b10000010011011011110100100100011101001111101000 :
(key == 11'b01010011010) ? 47'b10000010010010010111100100100011011100001101001 :
(key == 11'b01010011011) ? 47'b10000010001001010000110100100011001110011101111 :
(key == 11'b01010011100) ? 47'b10000010000000001010100100100011000000101111111 :
(key == 11'b01010011101) ? 47'b10000001110111000100110100100010110011000010111 :
(key == 11'b01010011110) ? 47'b10000001101101111111011100100010100101010110110 :
(key == 11'b01010011111) ? 47'b10000001100100111010011100100010010111101011100 :
(key == 11'b01010100000) ? 47'b10000001011011110101111100100010001010000001010 :
(key == 11'b01010100001) ? 47'b10000001010010110001110100100001111100011000000 :
(key == 11'b01010100010) ? 47'b10000001001001101110001100100001101110101111110 :
(key == 11'b01010100011) ? 47'b10000001000000101010111100100001100001001000100 :
(key == 11'b01010100100) ? 47'b10000000110111101000000100100001010011100010000 :
(key == 11'b01010100101) ? 47'b10000000101110100101101100100001000101111100101 :
(key == 11'b01010100110) ? 47'b10000000100101100011101100100000111000011000010 :
(key == 11'b01010100111) ? 47'b10000000011100100010001100100000101010110100110 :
(key == 11'b01010101000) ? 47'b10000000010011100001000100100000011101010010010 :
(key == 11'b01010101001) ? 47'b10000000001010100000010100100000001111110000101 :
(key == 11'b01010101010) ? 47'b10000000000001100000000100100000000010010000000 :
(key == 11'b01010101011) ? 47'b01111111111000100000001100011111110100110000010 :
(key == 11'b01010101100) ? 47'b01111111101111100000110100011111100111010001101 :
(key == 11'b01010101101) ? 47'b01111111100110100001110100011111011001110011111 :
(key == 11'b01010101110) ? 47'b01111111011101100011001100011111001100010111000 :
(key == 11'b01010101111) ? 47'b01111111010100100100111100011110111110111011000 :
(key == 11'b01010110000) ? 47'b01111111001011100111001100011110110001100000000 :
(key == 11'b01010110001) ? 47'b01111111000010101001111100011110100100000110001 :
(key == 11'b01010110010) ? 47'b01111110111001101100111100011110010110101101000 :
(key == 11'b01010110011) ? 47'b01111110110000110000011100011110001001010100111 :
(key == 11'b01010110100) ? 47'b01111110100111110100011100011101111011111101110 :
(key == 11'b01010110101) ? 47'b01111110011110111000101100011101101110100111011 :
(key == 11'b01010110110) ? 47'b01111110010101111101011100011101100001010010000 :
(key == 11'b01010110111) ? 47'b01111110001101000010101100011101010011111101110 :
(key == 11'b01010111000) ? 47'b01111110000100001000001100011101000110101010001 :
(key == 11'b01010111001) ? 47'b01111101111011001110001100011100111001010111101 :
(key == 11'b01010111010) ? 47'b01111101110010010100101100011100101100000110001 :
(key == 11'b01010111011) ? 47'b01111101101001011011011100011100011110110101011 :
(key == 11'b01010111100) ? 47'b01111101100000100010101100011100010001100101101 :
(key == 11'b01010111101) ? 47'b01111101010111101010010100011100000100010110110 :
(key == 11'b01010111110) ? 47'b01111101001110110010011100011011110111001000111 :
(key == 11'b01010111111) ? 47'b01111101000101111010111100011011101001111100000 :
(key == 11'b01011000000) ? 47'b01111100111101000011110100011011011100101111111 :
(key == 11'b01011000001) ? 47'b01111100110100001101001100011011001111100100110 :
(key == 11'b01011000010) ? 47'b01111100101011010110110100011011000010011010100 :
(key == 11'b01011000011) ? 47'b01111100100010100000111100011010110101010001001 :
(key == 11'b01011000100) ? 47'b01111100011001101011100100011010101000001000111 :
(key == 11'b01011000101) ? 47'b01111100010000110110011100011010011011000001010 :
(key == 11'b01011000110) ? 47'b01111100001000000001110100011010001101111010110 :
(key == 11'b01011000111) ? 47'b01111011111111001101100100011010000000110101000 :
(key == 11'b01011001000) ? 47'b01111011110110011001110100011001110011110000011 :
(key == 11'b01011001001) ? 47'b01111011101101100110010100011001100110101100100 :
(key == 11'b01011001010) ? 47'b01111011100100110011010100011001011001101001100 :
(key == 11'b01011001011) ? 47'b01111011011100000000110100011001001100100111101 :
(key == 11'b01011001100) ? 47'b01111011010011001110100100011000111111100110100 :
(key == 11'b01011001101) ? 47'b01111011001010011100110100011000110010100110010 :
(key == 11'b01011001110) ? 47'b01111011000001101011011100011000100101100111000 :
(key == 11'b01011001111) ? 47'b01111010111000111010011100011000011000101000100 :
(key == 11'b01011010000) ? 47'b01111010110000001001110100011000001011101010111 :
(key == 11'b01011010001) ? 47'b01111010100111011001101100010111111110101110011 :
(key == 11'b01011010010) ? 47'b01111010011110101001111100010111110001110010101 :
(key == 11'b01011010011) ? 47'b01111010010101111010100100010111100100110111111 :
(key == 11'b01011010100) ? 47'b01111010001101001011101100010111010111111110000 :
(key == 11'b01011010101) ? 47'b01111010000100011101000100010111001011000100111 :
(key == 11'b01011010110) ? 47'b01111001111011101110111100010110111110001100110 :
(key == 11'b01011010111) ? 47'b01111001110011000001001100010110110001010101100 :
(key == 11'b01011011000) ? 47'b01111001101010010011110100010110100100011111001 :
(key == 11'b01011011001) ? 47'b01111001100001100110111100010110010111101001110 :
(key == 11'b01011011010) ? 47'b01111001011000111010011100010110001010110101001 :
(key == 11'b01011011011) ? 47'b01111001010000001110001100010101111110000001011 :
(key == 11'b01011011100) ? 47'b01111001000111100010100100010101110001001110101 :
(key == 11'b01011011101) ? 47'b01111000111110110111001100010101100100011100101 :
(key == 11'b01011011110) ? 47'b01111000110110001100001100010101010111101011100 :
(key == 11'b01011011111) ? 47'b01111000101101100001101100010101001010111011011 :
(key == 11'b01011100000) ? 47'b01111000100100110111100100010100111110001100001 :
(key == 11'b01011100001) ? 47'b01111000011100001101110100010100110001011101110 :
(key == 11'b01011100010) ? 47'b01111000010011100100011100010100100100110000001 :
(key == 11'b01011100011) ? 47'b01111000001010111011100100010100011000000011101 :
(key == 11'b01011100100) ? 47'b01111000000010010010111100010100001011010111110 :
(key == 11'b01011100101) ? 47'b01110111111001101010110100010011111110101100111 :
(key == 11'b01011100110) ? 47'b01110111110001000011000100010011110010000010111 :
(key == 11'b01011100111) ? 47'b01110111101000011011101100010011100101011001101 :
(key == 11'b01011101000) ? 47'b01110111011111110100101100010011011000110001011 :
(key == 11'b01011101001) ? 47'b01110111010111001110000100010011001100001001110 :
(key == 11'b01011101010) ? 47'b01110111001110100111111100010010111111100011011 :
(key == 11'b01011101011) ? 47'b01110111000110000010001100010010110010111101101 :
(key == 11'b01011101100) ? 47'b01110110111101011100101100010010100110011000110 :
(key == 11'b01011101101) ? 47'b01110110110100110111101100010010011001110100110 :
(key == 11'b01011101110) ? 47'b01110110101100010011001100010010001101010001110 :
(key == 11'b01011101111) ? 47'b01110110100011101110111100010010000000101111100 :
(key == 11'b01011110000) ? 47'b01110110011011001011000100010001110100001110000 :
(key == 11'b01011110001) ? 47'b01110110010010100111101100010001100111101101101 :
(key == 11'b01011110010) ? 47'b01110110001010000100100100010001011011001101110 :
(key == 11'b01011110011) ? 47'b01110110000001100001111100010001001110101111000 :
(key == 11'b01011110100) ? 47'b01110101111000111111101100010001000010010001000 :
(key == 11'b01011110101) ? 47'b01110101110000011101110100010000110101110011111 :
(key == 11'b01011110110) ? 47'b01110101100111111100010100010000101001010111101 :
(key == 11'b01011110111) ? 47'b01110101011111011011001100010000011100111100010 :
(key == 11'b01011111000) ? 47'b01110101010110111010100100010000010000100001110 :
(key == 11'b01011111001) ? 47'b01110101001110011010001100010000000100001000000 :
(key == 11'b01011111010) ? 47'b01110101000101111010010100001111110111101111010 :
(key == 11'b01011111011) ? 47'b01110100111101011010101100001111101011010111000 :
(key == 11'b01011111100) ? 47'b01110100110100111011100100001111011110111111111 :
(key == 11'b01011111101) ? 47'b01110100101100011100110100001111010010101001101 :
(key == 11'b01011111110) ? 47'b01110100100011111110011100001111000110010100001 :
(key == 11'b01011111111) ? 47'b01110100011011100000011100001110111001111111100 :
(key == 11'b01100000000) ? 47'b01110100010011000010110100001110101101101011110 :
(key == 11'b01100000001) ? 47'b01110100001010100101100100001110100001011000110 :
(key == 11'b01100000010) ? 47'b01110100000010001000101100001110010101000110100 :
(key == 11'b01100000011) ? 47'b01110011111001101100001100001110001000110101010 :
(key == 11'b01100000100) ? 47'b01110011110001010000000100001101111100100100101 :
(key == 11'b01100000101) ? 47'b01110011101000110100011100001101110000010101001 :
(key == 11'b01100000110) ? 47'b01110011100000011001000100001101100100000110010 :
(key == 11'b01100000111) ? 47'b01110011010111111110001100001101010111111000011 :
(key == 11'b01100001000) ? 47'b01110011001111100011100100001101001011101011001 :
(key == 11'b01100001001) ? 47'b01110011000111001001011100001100111111011110111 :
(key == 11'b01100001010) ? 47'b01110010111110101111101100001100110011010011100 :
(key == 11'b01100001011) ? 47'b01110010110110010110001100001100100111001000110 :
(key == 11'b01100001100) ? 47'b01110010101101111101001100001100011010111111000 :
(key == 11'b01100001101) ? 47'b01110010100101100100100100001100001110110110000 :
(key == 11'b01100001110) ? 47'b01110010011101001100010100001100000010101101111 :
(key == 11'b01100001111) ? 47'b01110010010100110100010100001011110110100110011 :
(key == 11'b01100010000) ? 47'b01110010001100011100110100001011101010011111111 :
(key == 11'b01100010001) ? 47'b01110010000100000101101100001011011110011010001 :
(key == 11'b01100010010) ? 47'b01110001111011101110111100001011010010010101010 :
(key == 11'b01100010011) ? 47'b01110001110011011000100100001011000110010001010 :
(key == 11'b01100010100) ? 47'b01110001101011000010100100001010111010001110000 :
(key == 11'b01100010101) ? 47'b01110001100010101100111100001010101110001011100 :
(key == 11'b01100010110) ? 47'b01110001011010010111101100001010100010001001111 :
(key == 11'b01100010111) ? 47'b01110001010010000010110100001010010110001001001 :
(key == 11'b01100011000) ? 47'b01110001001001101110010100001010001010001001001 :
(key == 11'b01100011001) ? 47'b01110001000001011010001100001001111110001001111 :
(key == 11'b01100011010) ? 47'b01110000111001000110011100001001110010001011100 :
(key == 11'b01100011011) ? 47'b01110000110000110011000100001001100110001110000 :
(key == 11'b01100011100) ? 47'b01110000101000100000000100001001011010010001010 :
(key == 11'b01100011101) ? 47'b01110000100000001101011100001001001110010101010 :
(key == 11'b01100011110) ? 47'b01110000010111111011000100001001000010011001111 :
(key == 11'b01100011111) ? 47'b01110000001111101001001100001000110110011111101 :
(key == 11'b01100100000) ? 47'b01110000000111010111101100001000101010100110001 :
(key == 11'b01100100001) ? 47'b01101111111111000110100100001000011110101101011 :
(key == 11'b01100100010) ? 47'b01101111110110110101110100001000010010110101011 :
(key == 11'b01100100011) ? 47'b01101111101110100101011100001000000110111110011 :
(key == 11'b01100100100) ? 47'b01101111100110010101010100000111111011000111111 :
(key == 11'b01100100101) ? 47'b01101111011110000101101100000111101111010010011 :
(key == 11'b01100100110) ? 47'b01101111010101110110011100000111100011011101101 :
(key == 11'b01100100111) ? 47'b01101111001101100111011100000111010111101001100 :
(key == 11'b01100101000) ? 47'b01101111000101011000111100000111001011110110100 :
(key == 11'b01100101001) ? 47'b01101110111101001010101100000111000000000100000 :
(key == 11'b01100101010) ? 47'b01101110110100111100111100000110110100010010100 :
(key == 11'b01100101011) ? 47'b01101110101100101111011100000110101000100001101 :
(key == 11'b01100101100) ? 47'b01101110100100100010011100000110011100110001110 :
(key == 11'b01100101101) ? 47'b01101110011100010101101100000110010001000010100 :
(key == 11'b01100101110) ? 47'b01101110010100001001010100000110000101010100000 :
(key == 11'b01100101111) ? 47'b01101110001011111101010100000101111001100110011 :
(key == 11'b01100110000) ? 47'b01101110000011110001101100000101101101111001100 :
(key == 11'b01100110001) ? 47'b01101101111011100110011100000101100010001101011 :
(key == 11'b01100110010) ? 47'b01101101110011011011100100000101010110100010001 :
(key == 11'b01100110011) ? 47'b01101101101011010001000100000101001010110111101 :
(key == 11'b01100110100) ? 47'b01101101100011000110111100000100111111001110000 :
(key == 11'b01100110101) ? 47'b01101101011010111101000100000100110011100100111 :
(key == 11'b01100110110) ? 47'b01101101010010110011101100000100100111111100110 :
(key == 11'b01100110111) ? 47'b01101101001010101010100100000100011100010101011 :
(key == 11'b01100111000) ? 47'b01101101000010100001111100000100010000101110110 :
(key == 11'b01100111001) ? 47'b01101100111010011001100100000100000101001000111 :
(key == 11'b01100111010) ? 47'b01101100110010010001100100000011111001100011111 :
(key == 11'b01100111011) ? 47'b01101100101010001001111100000011101101111111100 :
(key == 11'b01100111100) ? 47'b01101100100010000010101100000011100010011100000 :
(key == 11'b01100111101) ? 47'b01101100011001111011110100000011010110111001010 :
(key == 11'b01100111110) ? 47'b01101100010001110101010100000011001011010111011 :
(key == 11'b01100111111) ? 47'b01101100001001101111000100000010111111110110000 :
(key == 11'b01101000000) ? 47'b01101100000001101001010100000010110100010101101 :
(key == 11'b01101000001) ? 47'b01101011111001100011110100000010101000110101111 :
(key == 11'b01101000010) ? 47'b01101011110001011110101100000010011101010111000 :
(key == 11'b01101000011) ? 47'b01101011101001011001111100000010010001111000110 :
(key == 11'b01101000100) ? 47'b01101011100001010101100100000010000110011011011 :
(key == 11'b01101000101) ? 47'b01101011011001010001100100000001111010111110110 :
(key == 11'b01101000110) ? 47'b01101011010001001101111100000001101111100011000 :
(key == 11'b01101000111) ? 47'b01101011001001001010100100000001100100000111110 :
(key == 11'b01101001000) ? 47'b01101011000001000111101100000001011000101101101 :
(key == 11'b01101001001) ? 47'b01101010111001000101000100000001001101010011111 :
(key == 11'b01101001010) ? 47'b01101010110001000010110100000001000001111011001 :
(key == 11'b01101001011) ? 47'b01101010101001000000111100000000110110100011000 :
(key == 11'b01101001100) ? 47'b01101010100000111111011100000000101011001011110 :
(key == 11'b01101001101) ? 47'b01101010011000111110010100000000011111110101010 :
(key == 11'b01101001110) ? 47'b01101010010000111101011100000000010100011111011 :
(key == 11'b01101001111) ? 47'b01101010001000111100111100000000001001001010010 :
(key == 11'b01101010000) ? 47'b01101010000000111100110011111111111101110101111 :
(key == 11'b01101010001) ? 47'b01101001111000111101000011111111110010100010011 :
(key == 11'b01101010010) ? 47'b01101001110000111101101011111111100111001111100 :
(key == 11'b01101010011) ? 47'b01101001101000111110101011111111011011111101100 :
(key == 11'b01101010100) ? 47'b01101001100000111111111011111111010000101100001 :
(key == 11'b01101010101) ? 47'b01101001011001000001100011111111000101011011100 :
(key == 11'b01101010110) ? 47'b01101001010001000011100011111110111010001011110 :
(key == 11'b01101010111) ? 47'b01101001001001000101111011111110101110111100101 :
(key == 11'b01101011000) ? 47'b01101001000001001000101011111110100011101110011 :
(key == 11'b01101011001) ? 47'b01101000111001001011101011111110011000100000110 :
(key == 11'b01101011010) ? 47'b01101000110001001111001011111110001101010100000 :
(key == 11'b01101011011) ? 47'b01101000101001010010111011111110000010000111111 :
(key == 11'b01101011100) ? 47'b01101000100001010111000011111101110110111100100 :
(key == 11'b01101011101) ? 47'b01101000011001011011011011111101101011110001110 :
(key == 11'b01101011110) ? 47'b01101000010001100000010011111101100000100111111 :
(key == 11'b01101011111) ? 47'b01101000001001100101011011111101010101011110110 :
(key == 11'b01101100000) ? 47'b01101000000001101010111011111101001010010110010 :
(key == 11'b01101100001) ? 47'b01100111111001110000110011111100111111001110101 :
(key == 11'b01101100010) ? 47'b01100111110001110110111011111100110100000111100 :
(key == 11'b01101100011) ? 47'b01100111101001111101100011111100101001000001011 :
(key == 11'b01101100100) ? 47'b01100111100010000100011011111100011101111011111 :
(key == 11'b01101100101) ? 47'b01100111011010001011101011111100010010110111001 :
(key == 11'b01101100110) ? 47'b01100111010010010011010011111100000111110011001 :
(key == 11'b01101100111) ? 47'b01100111001010011011001011111011111100101111110 :
(key == 11'b01101101000) ? 47'b01100111000010100011011011111011110001101101001 :
(key == 11'b01101101001) ? 47'b01100110111010101100000011111011100110101011010 :
(key == 11'b01101101010) ? 47'b01100110110010110101000011111011011011101010001 :
(key == 11'b01101101011) ? 47'b01100110101010111110010011111011010000101001101 :
(key == 11'b01101101100) ? 47'b01100110100011000111111011111011000101101001111 :
(key == 11'b01101101101) ? 47'b01100110011011010001111011111010111010101010111 :
(key == 11'b01101101110) ? 47'b01100110010011011100010011111010101111101100110 :
(key == 11'b01101101111) ? 47'b01100110001011100111000011111010100100101111010 :
(key == 11'b01101110000) ? 47'b01100110000011110010000011111010011001110010011 :
(key == 11'b01101110001) ? 47'b01100101111011111101011011111010001110110110011 :
(key == 11'b01101110010) ? 47'b01100101110100001001000011111010000011111010111 :
(key == 11'b01101110011) ? 47'b01100101101100010101001011111001111001000000010 :
(key == 11'b01101110100) ? 47'b01100101100100100001100011111001101110000110010 :
(key == 11'b01101110101) ? 47'b01100101011100101110010011111001100011001101001 :
(key == 11'b01101110110) ? 47'b01100101010100111011010011111001011000010100100 :
(key == 11'b01101110111) ? 47'b01100101001101001000110011111001001101011100110 :
(key == 11'b01101111000) ? 47'b01100101000101010110100011111001000010100101101 :
(key == 11'b01101111001) ? 47'b01100100111101100100100011111000110111101111001 :
(key == 11'b01101111010) ? 47'b01100100110101110011000011111000101100111001100 :
(key == 11'b01101111011) ? 47'b01100100101110000001110011111000100010000100100 :
(key == 11'b01101111100) ? 47'b01100100100110010000111011111000010111010000010 :
(key == 11'b01101111101) ? 47'b01100100011110100000010011111000001100011100101 :
(key == 11'b01101111110) ? 47'b01100100010110110000000011111000000001101001110 :
(key == 11'b01101111111) ? 47'b01100100001111000000001011110111110110110111101 :
(key == 11'b01110000000) ? 47'b01100100000111010000101011110111101100000110010 :
(key == 11'b01110000001) ? 47'b01100011111111100001011011110111100001010101011 :
(key == 11'b01110000010) ? 47'b01100011110111110010100011110111010110100101011 :
(key == 11'b01110000011) ? 47'b01100011110000000100000011110111001011110110000 :
(key == 11'b01110000100) ? 47'b01100011101000010101110011110111000001000111010 :
(key == 11'b01110000101) ? 47'b01100011100000100111111011110110110110011001011 :
(key == 11'b01110000110) ? 47'b01100011011000111010011011110110101011101100001 :
(key == 11'b01110000111) ? 47'b01100011010001001101010011110110100000111111101 :
(key == 11'b01110001000) ? 47'b01100011001001100000011011110110010110010011110 :
(key == 11'b01110001001) ? 47'b01100011000001110011110011110110001011101000100 :
(key == 11'b01110001010) ? 47'b01100010111010000111101011110110000000111110001 :
(key == 11'b01110001011) ? 47'b01100010110010011011110011110101110110010100010 :
(key == 11'b01110001100) ? 47'b01100010101010110000010011110101101011101011010 :
(key == 11'b01110001101) ? 47'b01100010100011000101000011110101100001000010110 :
(key == 11'b01110001110) ? 47'b01100010011011011010001011110101010110011011000 :
(key == 11'b01110001111) ? 47'b01100010010011101111101011110101001011110100001 :
(key == 11'b01110010000) ? 47'b01100010001100000101011011110101000001001101101 :
(key == 11'b01110010001) ? 47'b01100010000100011011100011110100110110101000000 :
(key == 11'b01110010010) ? 47'b01100001111100110010000011110100101100000011001 :
(key == 11'b01110010011) ? 47'b01100001110101001000110011110100100001011110110 :
(key == 11'b01110010100) ? 47'b01100001101101011111111011110100010110111011010 :
(key == 11'b01110010101) ? 47'b01100001100101110111011011110100001100011000011 :
(key == 11'b01110010110) ? 47'b01100001011110001111001011110100000001110110001 :
(key == 11'b01110010111) ? 47'b01100001010110100111010011110011110111010100101 :
(key == 11'b01110011000) ? 47'b01100001001110111111101011110011101100110011101 :
(key == 11'b01110011001) ? 47'b01100001000111011000011011110011100010010011011 :
(key == 11'b01110011010) ? 47'b01100000111111110001100011110011010111110100000 :
(key == 11'b01110011011) ? 47'b01100000111000001011000011110011001101010101010 :
(key == 11'b01110011100) ? 47'b01100000110000100100110011110011000010110111001 :
(key == 11'b01110011101) ? 47'b01100000101000111110110011110010111000011001100 :
(key == 11'b01110011110) ? 47'b01100000100001011001001011110010101101111100110 :
(key == 11'b01110011111) ? 47'b01100000011001110011111011110010100011100000101 :
(key == 11'b01110100000) ? 47'b01100000010010001111000011110010011001000101010 :
(key == 11'b01110100001) ? 47'b01100000001010101010011011110010001110101010100 :
(key == 11'b01110100010) ? 47'b01100000000011000110000011110010000100010000010 :
(key == 11'b01110100011) ? 47'b01011111111011100010000011110001111001110110110 :
(key == 11'b01110100100) ? 47'b01011111110011111110011011110001101111011110000 :
(key == 11'b01110100101) ? 47'b01011111101100011011001011110001100101000110000 :
(key == 11'b01110100110) ? 47'b01011111100100111000001011110001011010101110101 :
(key == 11'b01110100111) ? 47'b01011111011101010101011011110001010000010111110 :
(key == 11'b01110101000) ? 47'b01011111010101110011001011110001000110000001110 :
(key == 11'b01110101001) ? 47'b01011111001110010001000011110000111011101100001 :
(key == 11'b01110101010) ? 47'b01011111000110101111011011110000110001010111100 :
(key == 11'b01110101011) ? 47'b01011110111111001110000011110000100111000011011 :
(key == 11'b01110101100) ? 47'b01011110110111101100111011110000011100101111111 :
(key == 11'b01110101101) ? 47'b01011110110000001100001011110000010010011101001 :
(key == 11'b01110101110) ? 47'b01011110101000101011110011110000001000001011000 :
(key == 11'b01110101111) ? 47'b01011110100001001011101011101111111101111001100 :
(key == 11'b01110110000) ? 47'b01011110011001101011111011101111110011101000110 :
(key == 11'b01110110001) ? 47'b01011110010010001100011011101111101001011000100 :
(key == 11'b01110110010) ? 47'b01011110001010101101010011101111011111001001000 :
(key == 11'b01110110011) ? 47'b01011110000011001110100011101111010100111010011 :
(key == 11'b01110110100) ? 47'b01011101111011110000000011101111001010101100001 :
(key == 11'b01110110101) ? 47'b01011101110100010001110011101111000000011110100 :
(key == 11'b01110110110) ? 47'b01011101101100110100000011101110110110010001110 :
(key == 11'b01110110111) ? 47'b01011101100101010110011011101110101100000101100 :
(key == 11'b01110111000) ? 47'b01011101011101111001010011101110100001111010000 :
(key == 11'b01110111001) ? 47'b01011101010110011100010011101110010111101111000 :
(key == 11'b01110111010) ? 47'b01011101001110111111110011101110001101100100111 :
(key == 11'b01110111011) ? 47'b01011101000111100011100011101110000011011011010 :
(key == 11'b01110111100) ? 47'b01011101000000000111100011101101111001010010010 :
(key == 11'b01110111101) ? 47'b01011100111000101011111011101101101111001001111 :
(key == 11'b01110111110) ? 47'b01011100110001010000100011101101100101000010001 :
(key == 11'b01110111111) ? 47'b01011100101001110101100011101101011010111011001 :
(key == 11'b01111000000) ? 47'b01011100100010011010111011101101010000110100111 :
(key == 11'b01111000001) ? 47'b01011100011011000000100011101101000110101111001 :
(key == 11'b01111000010) ? 47'b01011100010011100110100011101100111100101010000 :
(key == 11'b01111000011) ? 47'b01011100001100001100110011101100110010100101101 :
(key == 11'b01111000100) ? 47'b01011100000100110011010011101100101000100001101 :
(key == 11'b01111000101) ? 47'b01011011111101011010001011101100011110011110100 :
(key == 11'b01111000110) ? 47'b01011011110110000001011011101100010100011100000 :
(key == 11'b01111000111) ? 47'b01011011101110101000111011101100001010011010001 :
(key == 11'b01111001000) ? 47'b01011011100111010000110011101100000000011000111 :
(key == 11'b01111001001) ? 47'b01011011011111111000111011101011110110011000010 :
(key == 11'b01111001010) ? 47'b01011011011000100001011011101011101100011000011 :
(key == 11'b01111001011) ? 47'b01011011010001001010001011101011100010011001000 :
(key == 11'b01111001100) ? 47'b01011011001001110011001011101011011000011010010 :
(key == 11'b01111001101) ? 47'b01011011000010011100101011101011001110011100010 :
(key == 11'b01111001110) ? 47'b01011010111011000110010011101011000100011110110 :
(key == 11'b01111001111) ? 47'b01011010110011110000010011101010111010100001111 :
(key == 11'b01111010000) ? 47'b01011010101100011010101011101010110000100101110 :
(key == 11'b01111010001) ? 47'b01011010100101000101010011101010100110101010010 :
(key == 11'b01111010010) ? 47'b01011010011101110000010011101010011100101111011 :
(key == 11'b01111010011) ? 47'b01011010010110011011100011101010010010110101001 :
(key == 11'b01111010100) ? 47'b01011010001111000111000011101010001000111011011 :
(key == 11'b01111010101) ? 47'b01011010000111110010111011101001111111000010011 :
(key == 11'b01111010110) ? 47'b01011010000000011111001011101001110101001010000 :
(key == 11'b01111010111) ? 47'b01011001111001001011101011101001101011010010010 :
(key == 11'b01111011000) ? 47'b01011001110001111000011011101001100001011011000 :
(key == 11'b01111011001) ? 47'b01011001101010100101100011101001010111100100100 :
(key == 11'b01111011010) ? 47'b01011001100011010010111011101001001101101110101 :
(key == 11'b01111011011) ? 47'b01011001011100000000101011101001000011111001011 :
(key == 11'b01111011100) ? 47'b01011001010100101110101011101000111010000100101 :
(key == 11'b01111011101) ? 47'b01011001001101011101000011101000110000010000101 :
(key == 11'b01111011110) ? 47'b01011001000110001011101011101000100110011101010 :
(key == 11'b01111011111) ? 47'b01011000111110111010101011101000011100101010100 :
(key == 11'b01111100000) ? 47'b01011000110111101001111011101000010010111000010 :
(key == 11'b01111100001) ? 47'b01011000110000011001011011101000001001000110101 :
(key == 11'b01111100010) ? 47'b01011000101001001001010011100111111111010101110 :
(key == 11'b01111100011) ? 47'b01011000100001111001100011100111110101100101100 :
(key == 11'b01111100100) ? 47'b01011000011010101010000011100111101011110101110 :
(key == 11'b01111100101) ? 47'b01011000010011011010110011100111100010000110101 :
(key == 11'b01111100110) ? 47'b01011000001100001011110011100111011000011000000 :
(key == 11'b01111100111) ? 47'b01011000000100111101010011100111001110101010011 :
(key == 11'b01111101000) ? 47'b01010111111101101110111011100111000100111101000 :
(key == 11'b01111101001) ? 47'b01010111110110100000111011100110111011010000011 :
(key == 11'b01111101010) ? 47'b01010111101111010011001011100110110001100100010 :
(key == 11'b01111101011) ? 47'b01010111101000000101110011100110100111111000110 :
(key == 11'b01111101100) ? 47'b01010111100000111000110011100110011110001110001 :
(key == 11'b01111101101) ? 47'b01010111011001101011111011100110010100100011110 :
(key == 11'b01111101110) ? 47'b01010111010010011111011011100110001010111010001 :
(key == 11'b01111101111) ? 47'b01010111001011010011010011100110000001010001010 :
(key == 11'b01111110000) ? 47'b01010111000100000111011011100101110111101000111 :
(key == 11'b01111110001) ? 47'b01010110111100111011110011100101101110000001000 :
(key == 11'b01111110010) ? 47'b01010110110101110000100011100101100100011001111 :
(key == 11'b01111110011) ? 47'b01010110101110100101100011100101011010110011010 :
(key == 11'b01111110100) ? 47'b01010110100111011010110011100101010001001101010 :
(key == 11'b01111110101) ? 47'b01010110100000010000011011100101000111100111111 :
(key == 11'b01111110110) ? 47'b01010110011001000110010011100100111110000011000 :
(key == 11'b01111110111) ? 47'b01010110010001111100100011100100110100011110111 :
(key == 11'b01111111000) ? 47'b01010110001010110011000011100100101010111011011 :
(key == 11'b01111111001) ? 47'b01010110000011101001111011100100100001011000011 :
(key == 11'b01111111010) ? 47'b01010101111100100000111011100100010111110101111 :
(key == 11'b01111111011) ? 47'b01010101110101011000011011100100001110010100010 :
(key == 11'b01111111100) ? 47'b01010101101110010000000011100100000100110011000 :
(key == 11'b01111111101) ? 47'b01010101100111001000000011100011111011010010011 :
(key == 11'b01111111110) ? 47'b01010101100000000000011011100011110001110010100 :
(key == 11'b01111111111) ? 47'b01010101011000111000111011100011101000010011000 :
(key == 11'b10000000000) ? 47'b01010101010001110001111011100011011110110100010 :
(key == 11'b10000000001) ? 47'b01010101001010101011000011100011010101010110000 :
(key == 11'b10000000010) ? 47'b01010101000011100100100011100011001011111000011 :
(key == 11'b10000000011) ? 47'b01010100111100011110010011100011000010011011010 :
(key == 11'b10000000100) ? 47'b01010100110101011000011011100010111000111110111 :
(key == 11'b10000000101) ? 47'b01010100101110010010110011100010101111100011000 :
(key == 11'b10000000110) ? 47'b01010100100111001101011011100010100110000111110 :
(key == 11'b10000000111) ? 47'b01010100100000001000011011100010011100101101001 :
(key == 11'b10000001000) ? 47'b01010100011001000011101011100010010011010011000 :
(key == 11'b10000001001) ? 47'b01010100010001111111001011100010001001111001100 :
(key == 11'b10000001010) ? 47'b01010100001010111011000011100010000000100000100 :
(key == 11'b10000001011) ? 47'b01010100000011110111001011100001110111001000010 :
(key == 11'b10000001100) ? 47'b01010011111100110011100011100001101101110000011 :
(key == 11'b10000001101) ? 47'b01010011110101110000010011100001100100011001010 :
(key == 11'b10000001110) ? 47'b01010011101110101101010011100001011011000010101 :
(key == 11'b10000001111) ? 47'b01010011100111101010100011100001010001101100101 :
(key == 11'b10000010000) ? 47'b01010011100000101000001011100001001000010111001 :
(key == 11'b10000010001) ? 47'b01010011011001100110000011100000111111000010011 :
(key == 11'b10000010010) ? 47'b01010011010010100100001011100000110101101110000 :
(key == 11'b10000010011) ? 47'b01010011001011100010101011100000101100011010011 :
(key == 11'b10000010100) ? 47'b01010011000100100001011011100000100011000111010 :
(key == 11'b10000010101) ? 47'b01010010111101100000100011100000011001110100110 :
(key == 11'b10000010110) ? 47'b01010010110110011111110011100000010000100010110 :
(key == 11'b10000010111) ? 47'b01010010101111011111011011100000000111010001010 :
(key == 11'b10000011000) ? 47'b01010010101000011111011011011111111110000000101 :
(key == 11'b10000011001) ? 47'b01010010100001011111100011011111110100110000010 :
(key == 11'b10000011010) ? 47'b01010010011010100000000011011111101011100000101 :
(key == 11'b10000011011) ? 47'b01010010010011100000111011011111100010010001101 :
(key == 11'b10000011100) ? 47'b01010010001100100001111011011111011001000011000 :
(key == 11'b10000011101) ? 47'b01010010000101100011010011011111001111110101001 :
(key == 11'b10000011110) ? 47'b01010001111110100100111011011111000110100111101 :
(key == 11'b10000011111) ? 47'b01010001110111100110111011011110111101011010111 :
(key == 11'b10000100000) ? 47'b01010001110000101001001011011110110100001110110 :
(key == 11'b10000100001) ? 47'b01010001101001101011101011011110101011000011000 :
(key == 11'b10000100010) ? 47'b01010001100010101110011011011110100001110111111 :
(key == 11'b10000100011) ? 47'b01010001011011110001100011011110011000101101011 :
(key == 11'b10000100100) ? 47'b01010001010100110100111011011110001111100011011 :
(key == 11'b10000100101) ? 47'b01010001001101111000100011011110000110011010000 :
(key == 11'b10000100110) ? 47'b01010001000110111100011011011101111101010001000 :
(key == 11'b10000100111) ? 47'b01010001000000000000101011011101110100001000110 :
(key == 11'b10000101000) ? 47'b01010000111001000101001011011101101011000001000 :
(key == 11'b10000101001) ? 47'b01010000110010001010000011011101100001111010000 :
(key == 11'b10000101010) ? 47'b01010000101011001111000011011101011000110011010 :
(key == 11'b10000101011) ? 47'b01010000100100010100011011011101001111101101010 :
(key == 11'b10000101100) ? 47'b01010000011101011010001011011101000110101000000 :
(key == 11'b10000101101) ? 47'b01010000010110100000000011011100111101100011000 :
(key == 11'b10000101110) ? 47'b01010000001111100110010011011100110100011110101 :
(key == 11'b10000101111) ? 47'b01010000001000101100110011011100101011011010111 :
(key == 11'b10000110000) ? 47'b01010000000001110011100011011100100010010111101 :
(key == 11'b10000110001) ? 47'b01001111111010111010101011011100011001010101000 :
(key == 11'b10000110010) ? 47'b01001111110100000001111011011100010000010010110 :
(key == 11'b10000110011) ? 47'b01001111101101001001100011011100000111010001001 :
(key == 11'b10000110100) ? 47'b01001111100110010001100011011011111110010000010 :
(key == 11'b10000110101) ? 47'b01001111011111011001101011011011110101001111101 :
(key == 11'b10000110110) ? 47'b01001111011000100010001011011011101100001111110 :
(key == 11'b10000110111) ? 47'b01001111010001101010111011011011100011010000011 :
(key == 11'b10000111000) ? 47'b01001111001010110100000011011011011010010001110 :
(key == 11'b10000111001) ? 47'b01001111000011111101010011011011010001010011011 :
(key == 11'b10000111010) ? 47'b01001110111101000110111011011011001000010101110 :
(key == 11'b10000111011) ? 47'b01001110110110010000110011011010111111011000101 :
(key == 11'b10000111100) ? 47'b01001110101111011010111011011010110110011011111 :
(key == 11'b10000111101) ? 47'b01001110101000100101011011011010101101100000000 :
(key == 11'b10000111110) ? 47'b01001110100001110000000011011010100100100100011 :
(key == 11'b10000111111) ? 47'b01001110011010111011000011011010011011101001011 :
(key == 11'b10001000000) ? 47'b01001110010100000110011011011010010010101111001 :
(key == 11'b10001000001) ? 47'b01001110001101010001111011011010001001110101001 :
(key == 11'b10001000010) ? 47'b01001110000110011101110011011010000000111011111 :
(key == 11'b10001000011) ? 47'b01001101111111101001111011011001111000000011001 :
(key == 11'b10001000100) ? 47'b01001101111000110110010011011001101111001010111 :
(key == 11'b10001000101) ? 47'b01001101110010000010111011011001100110010011001 :
(key == 11'b10001000110) ? 47'b01001101101011001111111011011001011101011100000 :
(key == 11'b10001000111) ? 47'b01001101100100011101000011011001010100100101010 :
(key == 11'b10001001000) ? 47'b01001101011101101010100011011001001011101111010 :
(key == 11'b10001001001) ? 47'b01001101010110111000010011011001000010111001101 :
(key == 11'b10001001010) ? 47'b01001101010000000110011011011000111010000100110 :
(key == 11'b10001001011) ? 47'b01001101001001010100101011011000110001010000010 :
(key == 11'b10001001100) ? 47'b01001101000010100011010011011000101000011100011 :
(key == 11'b10001001101) ? 47'b01001100111011110010001011011000011111101001000 :
(key == 11'b10001001110) ? 47'b01001100110101000001010011011000010110110110001 :
(key == 11'b10001001111) ? 47'b01001100101110010000110011011000001110000011111 :
(key == 11'b10001010000) ? 47'b01001100100111100000011011011000000101010010000 :
(key == 11'b10001010001) ? 47'b01001100100000110000011011010111111100100000110 :
(key == 11'b10001010010) ? 47'b01001100011010000000101011010111110011110000001 :
(key == 11'b10001010011) ? 47'b01001100010011010001001011010111101010111111111 :
(key == 11'b10001010100) ? 47'b01001100001100100010000011010111100010010000011 :
(key == 11'b10001010101) ? 47'b01001100000101110011000011010111011001100001001 :
(key == 11'b10001010110) ? 47'b01001011111111000100011011010111010000110010101 :
(key == 11'b10001010111) ? 47'b01001011111000010110000011010111001000000100101 :
(key == 11'b10001011000) ? 47'b01001011110001100111111011010110111111010111001 :
(key == 11'b10001011001) ? 47'b01001011101010111010000011010110110110101010000 :
(key == 11'b10001011010) ? 47'b01001011100100001100011011010110101101111101100 :
(key == 11'b10001011011) ? 47'b01001011011101011111001011010110100101010001101 :
(key == 11'b10001011100) ? 47'b01001011010110110010001011010110011100100110010 :
(key == 11'b10001011101) ? 47'b01001011010000000101011011010110010011111011011 :
(key == 11'b10001011110) ? 47'b01001011001001011000111011010110001011010001000 :
(key == 11'b10001011111) ? 47'b01001011000010101100101011010110000010100111001 :
(key == 11'b10001100000) ? 47'b01001010111100000000101011010101111001111101110 :
(key == 11'b10001100001) ? 47'b01001010110101010101000011010101110001010101001 :
(key == 11'b10001100010) ? 47'b01001010101110101001101011010101101000101100111 :
(key == 11'b10001100011) ? 47'b01001010100111111110100011010101100000000101001 :
(key == 11'b10001100100) ? 47'b01001010100001010011101011010101010111011101111 :
(key == 11'b10001100101) ? 47'b01001010011010101001000011010101001110110111010 :
(key == 11'b10001100110) ? 47'b01001010010011111110101011010101000110010001000 :
(key == 11'b10001100111) ? 47'b01001010001101010100101011010100111101101011011 :
(key == 11'b10001101000) ? 47'b01001010000110101010111011010100110101000110011 :
(key == 11'b10001101001) ? 47'b01001010000000000001010011010100101100100001101 :
(key == 11'b10001101010) ? 47'b01001001111001011000000011010100100011111101100 :
(key == 11'b10001101011) ? 47'b01001001110010101111000011010100011011011001111 :
(key == 11'b10001101100) ? 47'b01001001101100000110011011010100010010110111000 :
(key == 11'b10001101101) ? 47'b01001001100101011101111011010100001010010100011 :
(key == 11'b10001101110) ? 47'b01001001011110110101101011010100000001110010010 :
(key == 11'b10001101111) ? 47'b01001001011000001101110011010011111001010000110 :
(key == 11'b10001110000) ? 47'b01001001010001100110001011010011110000101111111 :
(key == 11'b10001110001) ? 47'b01001001001010111110110011010011101000001111011 :
(key == 11'b10001110010) ? 47'b01001001000100010111101011010011011111101111011 :
(key == 11'b10001110011) ? 47'b01001000111101110000110011010011010111001111111 :
(key == 11'b10001110100) ? 47'b01001000110111001010001011010011001110110000111 :
(key == 11'b10001110101) ? 47'b01001000110000100011110011010011000110010010011 :
(key == 11'b10001110110) ? 47'b01001000101001111101110011010010111101110100100 :
(key == 11'b10001110111) ? 47'b01001000100011010111111011010010110101010111000 :
(key == 11'b10001111000) ? 47'b01001000011100110010011011010010101100111010001 :
(key == 11'b10001111001) ? 47'b01001000010110001101001011010010100100011101110 :
(key == 11'b10001111010) ? 47'b01001000001111101000001011010010011100000001111 :
(key == 11'b10001111011) ? 47'b01001000001001000011011011010010010011100110100 :
(key == 11'b10001111100) ? 47'b01001000000010011110111011010010001011001011100 :
(key == 11'b10001111101) ? 47'b01000111111011111010101011010010000010110001001 :
(key == 11'b10001111110) ? 47'b01000111110101010110110011010001111010010111011 :
(key == 11'b10001111111) ? 47'b01000111101110110011000011010001110001111101111 :
(key == 11'b10010000000) ? 47'b01000111101000001111101011010001101001100101001 :
(key == 11'b10010000001) ? 47'b01000111100001101100011011010001100001001100101 :
(key == 11'b10010000010) ? 47'b01000111011011001001100011010001011000110100110 :
(key == 11'b10010000011) ? 47'b01000111010100100110111011010001010000011101100 :
(key == 11'b10010000100) ? 47'b01000111001110000100100011010001001000000110101 :
(key == 11'b10010000101) ? 47'b01000111000111100010011011010000111111110000010 :
(key == 11'b10010000110) ? 47'b01000111000001000000100011010000110111011010011 :
(key == 11'b10010000111) ? 47'b01000110111010011110111011010000101111000101000 :
(key == 11'b10010001000) ? 47'b01000110110011111101101011010000100110110000010 :
(key == 11'b10010001001) ? 47'b01000110101101011100100011010000011110011011110 :
(key == 11'b10010001010) ? 47'b01000110100110111011101011010000010110000111111 :
(key == 11'b10010001011) ? 47'b01000110100000011011001011010000001101110100101 :
(key == 11'b10010001100) ? 47'b01000110011001111010110011010000000101100001101 :
(key == 11'b10010001101) ? 47'b01000110010011011010110011001111111101001111010 :
(key == 11'b10010001110) ? 47'b01000110001100111011000011001111110100111101011 :
(key == 11'b10010001111) ? 47'b01000110000110011011100011001111101100101100001 :
(key == 11'b10010010000) ? 47'b01000101111111111100001011001111100100011011000 :
(key == 11'b10010010001) ? 47'b01000101111001011101001011001111011100001010101 :
(key == 11'b10010010010) ? 47'b01000101110010111110011011001111010011111010110 :
(key == 11'b10010010011) ? 47'b01000101101100011111111011001111001011101011010 :
(key == 11'b10010010100) ? 47'b01000101100110000001110011001111000011011100100 :
(key == 11'b10010010101) ? 47'b01000101011111100011110011001110111011001110000 :
(key == 11'b10010010110) ? 47'b01000101011001000110000011001110110011000000001 :
(key == 11'b10010010111) ? 47'b01000101010010101000100011001110101010110010101 :
(key == 11'b10010011000) ? 47'b01000101001100001011011011001110100010100101110 :
(key == 11'b10010011001) ? 47'b01000101000101101110011011001110011010011001001 :
(key == 11'b10010011010) ? 47'b01000100111111010001101011001110010010001101001 :
(key == 11'b10010011011) ? 47'b01000100111000110101010011001110001010000001101 :
(key == 11'b10010011100) ? 47'b01000100110010011001000011001110000001110110101 :
(key == 11'b10010011101) ? 47'b01000100101011111101001011001101111001101100001 :
(key == 11'b10010011110) ? 47'b01000100100101100001011011001101110001100010000 :
(key == 11'b10010011111) ? 47'b01000100011111000110000011001101101001011000100 :
(key == 11'b10010100000) ? 47'b01000100011000101010111011001101100001001111011 :
(key == 11'b10010100001) ? 47'b01000100010010001111111011001101011001000110110 :
(key == 11'b10010100010) ? 47'b01000100001011110101010011001101010000111110101 :
(key == 11'b10010100011) ? 47'b01000100000101011010111011001101001000110111000 :
(key == 11'b10010100100) ? 47'b01000011111111000000110011001101000000101111111 :
(key == 11'b10010100101) ? 47'b01000011111000100110111011001100111000101001010 :
(key == 11'b10010100110) ? 47'b01000011110010001101001011001100110000100011000 :
(key == 11'b10010100111) ? 47'b01000011101011110011110011001100101000011101010 :
(key == 11'b10010101000) ? 47'b01000011100101011010101011001100100000011000000 :
(key == 11'b10010101001) ? 47'b01000011011111000001110011001100011000010011010 :
(key == 11'b10010101010) ? 47'b01000011011000101001001011001100010000001111000 :
(key == 11'b10010101011) ? 47'b01000011010010010000110011001100001000001011010 :
(key == 11'b10010101100) ? 47'b01000011001011111000101011001100000000001000000 :
(key == 11'b10010101101) ? 47'b01000011000101100000110011001011111000000101001 :
(key == 11'b10010101110) ? 47'b01000010111111001001001011001011110000000010110 :
(key == 11'b10010101111) ? 47'b01000010111000110001110011001011101000000000111 :
(key == 11'b10010110000) ? 47'b01000010110010011010101011001011011111111111011 :
(key == 11'b10010110001) ? 47'b01000010101100000011110011001011010111111110100 :
(key == 11'b10010110010) ? 47'b01000010100101101101001011001011001111111110000 :
(key == 11'b10010110011) ? 47'b01000010011111010110110011001011000111111110000 :
(key == 11'b10010110100) ? 47'b01000010011001000000101011001010111111111110100 :
(key == 11'b10010110101) ? 47'b01000010010010101010110011001010110111111111011 :
(key == 11'b10010110110) ? 47'b01000010001100010101001011001010110000000000111 :
(key == 11'b10010110111) ? 47'b01000010000101111111110011001010101000000010110 :
(key == 11'b10010111000) ? 47'b01000001111111101010101011001010100000000101001 :
(key == 11'b10010111001) ? 47'b01000001111001010101110011001010011000000111111 :
(key == 11'b10010111010) ? 47'b01000001110011000001001011001010010000001011010 :
(key == 11'b10010111011) ? 47'b01000001101100101100110011001010001000001111000 :
(key == 11'b10010111100) ? 47'b01000001100110011000101011001010000000010011010 :
(key == 11'b10010111101) ? 47'b01000001100000000100110011001001111000010111111 :
(key == 11'b10010111110) ? 47'b01000001011001110001001011001001110000011101001 :
(key == 11'b10010111111) ? 47'b01000001010011011101101011001001101000100010101 :
(key == 11'b10011000000) ? 47'b01000001001101001010100011001001100000101000110 :
(key == 11'b10011000001) ? 47'b01000001000110110111101011001001011000101111010 :
(key == 11'b10011000010) ? 47'b01000001000000100101000011001001010000110110011 :
(key == 11'b10011000011) ? 47'b01000000111010010010101011001001001000111101111 :
(key == 11'b10011000100) ? 47'b01000000110100000000011011001001000001000101110 :
(key == 11'b10011000101) ? 47'b01000000101101101110100011001000111001001110001 :
(key == 11'b10011000110) ? 47'b01000000100111011100111011001000110001010111001 :
(key == 11'b10011000111) ? 47'b01000000100001001011011011001000101001100000011 :
(key == 11'b10011001000) ? 47'b01000000011010111010010011001000100001101010010 :
(key == 11'b10011001001) ? 47'b01000000010100101001011011001000011001110100100 :
(key == 11'b10011001010) ? 47'b01000000001110011000101011001000010001111111001 :
(key == 11'b10011001011) ? 47'b01000000001000001000010011001000001010001010011 :
(key == 11'b10011001100) ? 47'b01000000000001111000000011001000000010010110000 :
(key == 11'b10011001101) ? 47'b00111111111011101000000011000111111010100010000 :
(key == 11'b10011001110) ? 47'b00111111110101011000011011000111110010101110101 :
(key == 11'b10011001111) ? 47'b00111111101111001000111011000111101010111011101 :
(key == 11'b10011010000) ? 47'b00111111101000111001101011000111100011001001000 :
(key == 11'b10011010001) ? 47'b00111111100010101010110011000111011011010111001 :
(key == 11'b10011010010) ? 47'b00111111011100011100000011000111010011100101100 :
(key == 11'b10011010011) ? 47'b00111111010110001101100011000111001011110100010 :
(key == 11'b10011010100) ? 47'b00111111001111111111010011000111000100000011100 :
(key == 11'b10011010101) ? 47'b00111111001001110001010011000110111100010011010 :
(key == 11'b10011010110) ? 47'b00111111000011100011100011000110110100100011100 :
(key == 11'b10011010111) ? 47'b00111110111101010101111011000110101100110100000 :
(key == 11'b10011011000) ? 47'b00111110110111001000101011000110100101000101001 :
(key == 11'b10011011001) ? 47'b00111110110000111011101011000110011101010110110 :
(key == 11'b10011011010) ? 47'b00111110101010101110111011000110010101101000110 :
(key == 11'b10011011011) ? 47'b00111110100100100010010011000110001101111011001 :
(key == 11'b10011011100) ? 47'b00111110011110010110000011000110000110001110001 :
(key == 11'b10011011101) ? 47'b00111110011000001001111011000101111110100001011 :
(key == 11'b10011011110) ? 47'b00111110010001111110000011000101110110110101001 :
(key == 11'b10011011111) ? 47'b00111110001011110010100011000101101111001001100 :
(key == 11'b10011100000) ? 47'b00111110000101100111001011000101100111011110001 :
(key == 11'b10011100001) ? 47'b00111101111111011100000011000101011111110011010 :
(key == 11'b10011100010) ? 47'b00111101111001010001001011000101011000001000111 :
(key == 11'b10011100011) ? 47'b00111101110011000110100011000101010000011110111 :
(key == 11'b10011100100) ? 47'b00111101101100111100001011000101001000110101011 :
(key == 11'b10011100101) ? 47'b00111101100110110001111011000101000001001100001 :
(key == 11'b10011100110) ? 47'b00111101100000101000000011000100111001100011101 :
(key == 11'b10011100111) ? 47'b00111101011010011110011011000100110001111011100 :
(key == 11'b10011101000) ? 47'b00111101010100010100111011000100101010010011101 :
(key == 11'b10011101001) ? 47'b00111101001110001011101011000100100010101100010 :
(key == 11'b10011101010) ? 47'b00111101001000000010110011000100011011000101100 :
(key == 11'b10011101011) ? 47'b00111101000001111010000011000100010011011111000 :
(key == 11'b10011101100) ? 47'b00111100111011110001100011000100001011111001000 :
(key == 11'b10011101101) ? 47'b00111100110101101001010011000100000100010011100 :
(key == 11'b10011101110) ? 47'b00111100101111100001010011000011111100101110011 :
(key == 11'b10011101111) ? 47'b00111100101001011001100011000011110101001001110 :
(key == 11'b10011110000) ? 47'b00111100100011010001111011000011101101100101100 :
(key == 11'b10011110001) ? 47'b00111100011101001010101011000011100110000001110 :
(key == 11'b10011110010) ? 47'b00111100010111000011100011000011011110011110011 :
(key == 11'b10011110011) ? 47'b00111100010000111100110011000011010110111011100 :
(key == 11'b10011110100) ? 47'b00111100001010110110001011000011001111011001000 :
(key == 11'b10011110101) ? 47'b00111100000100101111110011000011000111110111000 :
(key == 11'b10011110110) ? 47'b00111011111110101001101011000011000000010101011 :
(key == 11'b10011110111) ? 47'b00111011111000100011110011000010111000110100010 :
(key == 11'b10011111000) ? 47'b00111011110010011110000011000010110001010011011 :
(key == 11'b10011111001) ? 47'b00111011101100011000101011000010101001110011001 :
(key == 11'b10011111010) ? 47'b00111011100110010011011011000010100010010011001 :
(key == 11'b10011111011) ? 47'b00111011100000001110100011000010011010110011111 :
(key == 11'b10011111100) ? 47'b00111011011010001001110011000010010011010100110 :
(key == 11'b10011111101) ? 47'b00111011010100000101010011000010001011110110010 :
(key == 11'b10011111110) ? 47'b00111011001110000001000011000010000100011000001 :
(key == 11'b10011111111) ? 47'b00111011000111111101000011000001111100111010011 :
(key == 11'b10100000000) ? 47'b00111011000001111001010011000001110101011101001 :
(key == 11'b10100000001) ? 47'b00111010111011110101101011000001101110000000010 :
(key == 11'b10100000010) ? 47'b00111010110101110010011011000001100110100011111 :
(key == 11'b10100000011) ? 47'b00111010101111101111010011000001011111000111111 :
(key == 11'b10100000100) ? 47'b00111010101001101100011011000001010111101100010 :
(key == 11'b10100000101) ? 47'b00111010100011101001110011000001010000010001001 :
(key == 11'b10100000110) ? 47'b00111010011101100111011011000001001000110110100 :
(key == 11'b10100000111) ? 47'b00111010010111100101010011000001000001011100010 :
(key == 11'b10100001000) ? 47'b00111010010001100011010011000000111010000010010 :
(key == 11'b10100001001) ? 47'b00111010001011100001101011000000110010101001000 :
(key == 11'b10100001010) ? 47'b00111010000101100000001011000000101011001111111 :
(key == 11'b10100001011) ? 47'b00111001111111011110111011000000100011110111011 :
(key == 11'b10100001100) ? 47'b00111001111001011101111011000000011100011111010 :
(key == 11'b10100001101) ? 47'b00111001110011011101001011000000010101000111100 :
(key == 11'b10100001110) ? 47'b00111001101101011100100011000000001101110000001 :
(key == 11'b10100001111) ? 47'b00111001100111011100010011000000000110011001010 :
(key == 11'b10100010000) ? 47'b00111001100001011100001010111111111111000010110 :
(key == 11'b10100010001) ? 47'b00111001011011011100010010111111110111101100110 :
(key == 11'b10100010010) ? 47'b00111001010101011100101010111111110000010111001 :
(key == 11'b10100010011) ? 47'b00111001001111011101010010111111101001000010000 :
(key == 11'b10100010100) ? 47'b00111001001001011110001010111111100001101101010 :
(key == 11'b10100010101) ? 47'b00111001000011011111001010111111011010011000110 :
(key == 11'b10100010110) ? 47'b00111000111101100000100010111111010011000101000 :
(key == 11'b10100010111) ? 47'b00111000110111100010000010111111001011110001011 :
(key == 11'b10100011000) ? 47'b00111000110001100011110010111111000100011110011 :
(key == 11'b10100011001) ? 47'b00111000101011100101110010111110111101001011110 :
(key == 11'b10100011010) ? 47'b00111000100101100111111010111110110101111001011 :
(key == 11'b10100011011) ? 47'b00111000011111101010011010111110101110100111101 :
(key == 11'b10100011100) ? 47'b00111000011001101101000010111110100111010110001 :
(key == 11'b10100011101) ? 47'b00111000010011101111111010111110100000000101001 :
(key == 11'b10100011110) ? 47'b00111000001101110011000010111110011000110100100 :
(key == 11'b10100011111) ? 47'b00111000000111110110011010111110010001100100011 :
(key == 11'b10100100000) ? 47'b00111000000001111001111010111110001010010100100 :
(key == 11'b10100100001) ? 47'b00110111111011111101101010111110000011000101001 :
(key == 11'b10100100010) ? 47'b00110111110110000001110010111101111011110110010 :
(key == 11'b10100100011) ? 47'b00110111110000000101111010111101110100100111101 :
(key == 11'b10100100100) ? 47'b00110111101010001010011010111101101101011001100 :
(key == 11'b10100100101) ? 47'b00110111100100001111001010111101100110001011111 :
(key == 11'b10100100110) ? 47'b00110111011110010100000010111101011110111110100 :
(key == 11'b10100100111) ? 47'b00110111011000011001001010111101010111110001101 :
(key == 11'b10100101000) ? 47'b00110111010010011110100010111101010000100101010 :
(key == 11'b10100101001) ? 47'b00110111001100100100001010111101001001011001001 :
(key == 11'b10100101010) ? 47'b00110111000110101010000010111101000010001101101 :
(key == 11'b10100101011) ? 47'b00110111000000110000000010111100111011000010010 :
(key == 11'b10100101100) ? 47'b00110110111010110110010010111100110011110111011 :
(key == 11'b10100101101) ? 47'b00110110110100111100110010111100101100101101000 :
(key == 11'b10100101110) ? 47'b00110110101111000011100010111100100101100011000 :
(key == 11'b10100101111) ? 47'b00110110101001001010011010111100011110011001011 :
(key == 11'b10100110000) ? 47'b00110110100011010001100010111100010111010000001 :
(key == 11'b10100110001) ? 47'b00110110011101011001000010111100010000000111011 :
(key == 11'b10100110010) ? 47'b00110110010111100000100010111100001000111110111 :
(key == 11'b10100110011) ? 47'b00110110010001101000011010111100000001110111000 :
(key == 11'b10100110100) ? 47'b00110110001011110000100010111011111010101111100 :
(key == 11'b10100110101) ? 47'b00110110000101111000110010111011110011101000010 :
(key == 11'b10100110110) ? 47'b00110110000000000001010010111011101100100001100 :
(key == 11'b10100110111) ? 47'b00110101111010001001111010111011100101011011000 :
(key == 11'b10100111000) ? 47'b00110101110100010010111010111011011110010101001 :
(key == 11'b10100111001) ? 47'b00110101101110011100000010111011010111001111100 :
(key == 11'b10100111010) ? 47'b00110101101000100101011010111011010000001010010 :
(key == 11'b10100111011) ? 47'b00110101100010101111000010111011001001000101100 :
(key == 11'b10100111100) ? 47'b00110101011100111000111010111011000010000001010 :
(key == 11'b10100111101) ? 47'b00110101010111000010111010111010111010111101010 :
(key == 11'b10100111110) ? 47'b00110101010001001101001010111010110011111001101 :
(key == 11'b10100111111) ? 47'b00110101001011010111101010111010101100110110100 :
(key == 11'b10101000000) ? 47'b00110101000101100010011010111010100101110011110 :
(key == 11'b10101000001) ? 47'b00110100111111101101010010111010011110110001011 :
(key == 11'b10101000010) ? 47'b00110100111001111000100010111010010111101111100 :
(key == 11'b10101000011) ? 47'b00110100110100000011110010111010010000101101110 :
(key == 11'b10101000100) ? 47'b00110100101110001111011010111010001001101100101 :
(key == 11'b10101000101) ? 47'b00110100101000011011010010111010000010101100000 :
(key == 11'b10101000110) ? 47'b00110100100010100111010010111001111011101011100 :
(key == 11'b10101000111) ? 47'b00110100011100110011100010111001110100101011100 :
(key == 11'b10101001000) ? 47'b00110100010110111111111010111001101101101011111 :
(key == 11'b10101001001) ? 47'b00110100010001001100101010111001100110101100110 :
(key == 11'b10101001010) ? 47'b00110100001011011001100010111001011111101101111 :
(key == 11'b10101001011) ? 47'b00110100000101100110101010111001011000101111100 :
(key == 11'b10101001100) ? 47'b00110011111111110100000010111001010001110001100 :
(key == 11'b10101001101) ? 47'b00110011111010000001100010111001001010110011111 :
(key == 11'b10101001110) ? 47'b00110011110100001111010010111001000011110110101 :
(key == 11'b10101001111) ? 47'b00110011101110011101010010111000111100111001110 :
(key == 11'b10101010000) ? 47'b00110011101000101011100010111000110101111101011 :
(key == 11'b10101010001) ? 47'b00110011100010111001111010111000101111000001010 :
(key == 11'b10101010010) ? 47'b00110011011101001000100010111000101000000101101 :
(key == 11'b10101010011) ? 47'b00110011010111010111011010111000100001001010011 :
(key == 11'b10101010100) ? 47'b00110011010001100110100010111000011010001111100 :
(key == 11'b10101010101) ? 47'b00110011001011110101110010111000010011010101000 :
(key == 11'b10101010110) ? 47'b00110011000110000101010010111000001100011010111 :
(key == 11'b10101010111) ? 47'b00110011000000010101000010111000000101100001001 :
(key == 11'b10101011000) ? 47'b00110010111010100100111010110111111110100111110 :
(key == 11'b10101011001) ? 47'b00110010110100110101001010110111110111101110111 :
(key == 11'b10101011010) ? 47'b00110010101111000101100010110111110000110110011 :
(key == 11'b10101011011) ? 47'b00110010101001010110000010110111101001111110001 :
(key == 11'b10101011100) ? 47'b00110010100011100110111010110111100011000110011 :
(key == 11'b10101011101) ? 47'b00110010011101110111111010110111011100001111000 :
(key == 11'b10101011110) ? 47'b00110010011000001001000010110111010101010111111 :
(key == 11'b10101011111) ? 47'b00110010010010011010100010110111001110100001010 :
(key == 11'b10101100000) ? 47'b00110010001100101100001010110111000111101011000 :
(key == 11'b10101100001) ? 47'b00110010000110111110000010110111000000110101001 :
(key == 11'b10101100010) ? 47'b00110010000001010000001010110110111001111111110 :
(key == 11'b10101100011) ? 47'b00110001111011100010011010110110110011001010101 :
(key == 11'b10101100100) ? 47'b00110001110101110100111010110110101100010101111 :
(key == 11'b10101100101) ? 47'b00110001110000000111101010110110100101100001101 :
(key == 11'b10101100110) ? 47'b00110001101010011010100010110110011110101101100 :
(key == 11'b10101100111) ? 47'b00110001100100101101110010110110010111111010001 :
(key == 11'b10101101000) ? 47'b00110001011111000001000010110110010001000110110 :
(key == 11'b10101101001) ? 47'b00110001011001010100101010110110001010010100000 :
(key == 11'b10101101010) ? 47'b00110001010011101000011010110110000011100001101 :
(key == 11'b10101101011) ? 47'b00110001001101111100011010110101111100101111100 :
(key == 11'b10101101100) ? 47'b00110001001000010000101010110101110101111101111 :
(key == 11'b10101101101) ? 47'b00110001000010100101000010110101101111001100101 :
(key == 11'b10101101110) ? 47'b00110000111100111001101010110101101000011011101 :
(key == 11'b10101101111) ? 47'b00110000110111001110100010110101100001101011001 :
(key == 11'b10101110000) ? 47'b00110000110001100011100010110101011010111010111 :
(key == 11'b10101110001) ? 47'b00110000101011111000111010110101010100001011010 :
(key == 11'b10101110010) ? 47'b00110000100110001110010010110101001101011011110 :
(key == 11'b10101110011) ? 47'b00110000100000100100000010110101000110101100110 :
(key == 11'b10101110100) ? 47'b00110000011010111001111010110100111111111110001 :
(key == 11'b10101110101) ? 47'b00110000010101010000000010110100111001001111111 :
(key == 11'b10101110110) ? 47'b00110000001111100110010010110100110010100001111 :
(key == 11'b10101110111) ? 47'b00110000001001111100111010110100101011110100100 :
(key == 11'b10101111000) ? 47'b00110000000100010011100010110100100101000111001 :
(key == 11'b10101111001) ? 47'b00101111111110101010100010110100011110011010100 :
(key == 11'b10101111010) ? 47'b00101111111001000001101010110100010111101110000 :
(key == 11'b10101111011) ? 47'b00101111110011011001000010110100010001000010000 :
(key == 11'b10101111100) ? 47'b00101111101101110000101010110100001010010110011 :
(key == 11'b10101111101) ? 47'b00101111101000001000011010110100000011101011000 :
(key == 11'b10101111110) ? 47'b00101111100010100000011010110011111101000000001 :
(key == 11'b10101111111) ? 47'b00101111011100111000101010110011110110010101101 :
(key == 11'b10110000000) ? 47'b00101111010111010001000010110011101111101011011 :
(key == 11'b10110000001) ? 47'b00101111010001101001101010110011101001000001101 :
(key == 11'b10110000010) ? 47'b00101111001100000010011010110011100010011000001 :
(key == 11'b10110000011) ? 47'b00101111000110011011011010110011011011101111000 :
(key == 11'b10110000100) ? 47'b00101111000000110100101010110011010101000110010 :
(key == 11'b10110000101) ? 47'b00101110111011001110001010110011001110011110000 :
(key == 11'b10110000110) ? 47'b00101110110101100111110010110011000111110110000 :
(key == 11'b10110000111) ? 47'b00101110110000000001101010110011000001001110011 :
(key == 11'b10110001000) ? 47'b00101110101010011011110010110010111010100111010 :
(key == 11'b10110001001) ? 47'b00101110100100110110000010110010110100000000011 :
(key == 11'b10110001010) ? 47'b00101110011111010000100010110010101101011001111 :
(key == 11'b10110001011) ? 47'b00101110011001101011001010110010100110110011101 :
(key == 11'b10110001100) ? 47'b00101110010100000110000010110010100000001101111 :
(key == 11'b10110001101) ? 47'b00101110001110100001001010110010011001101000100 :
(key == 11'b10110001110) ? 47'b00101110001000111100011010110010010011000011011 :
(key == 11'b10110001111) ? 47'b00101110000011010111111010110010001100011110101 :
(key == 11'b10110010000) ? 47'b00101101111101110011101010110010000101111010011 :
(key == 11'b10110010001) ? 47'b00101101111000001111100010110001111111010110011 :
(key == 11'b10110010010) ? 47'b00101101110010101011101010110001111000110010110 :
(key == 11'b10110010011) ? 47'b00101101101101001000000010110001110010001111101 :
(key == 11'b10110010100) ? 47'b00101101100111100100100010110001101011101100110 :
(key == 11'b10110010101) ? 47'b00101101100010000001010010110001100101001010010 :
(key == 11'b10110010110) ? 47'b00101101011100011110010010110001011110101000001 :
(key == 11'b10110010111) ? 47'b00101101010110111011011010110001011000000110010 :
(key == 11'b10110011000) ? 47'b00101101010001011000110010110001010001100100111 :
(key == 11'b10110011001) ? 47'b00101101001011110110010010110001001011000011110 :
(key == 11'b10110011010) ? 47'b00101101000110010100000010110001000100100011000 :
(key == 11'b10110011011) ? 47'b00101101000000110010000010110000111110000010110 :
(key == 11'b10110011100) ? 47'b00101100111011010000001010110000110111100010110 :
(key == 11'b10110011101) ? 47'b00101100110101101110100010110000110001000011001 :
(key == 11'b10110011110) ? 47'b00101100110000001101001010110000101010100011111 :
(key == 11'b10110011111) ? 47'b00101100101010101011111010110000100100000101000 :
(key == 11'b10110100000) ? 47'b00101100100101001010111010110000011101100110011 :
(key == 11'b10110100001) ? 47'b00101100011111101010000010110000010111001000001 :
(key == 11'b10110100010) ? 47'b00101100011010001001011010110000010000101010010 :
(key == 11'b10110100011) ? 47'b00101100010100101001000010110000001010001100111 :
(key == 11'b10110100100) ? 47'b00101100001111001000110010110000000011101111101 :
(key == 11'b10110100101) ? 47'b00101100001001101000110010101111111101010010111 :
(key == 11'b10110100110) ? 47'b00101100000100001000111010101111110110110110011 :
(key == 11'b10110100111) ? 47'b00101011111110101001010010101111110000011010010 :
(key == 11'b10110101000) ? 47'b00101011111001001001111010101111101001111110101 :
(key == 11'b10110101001) ? 47'b00101011110011101010101010101111100011100011010 :
(key == 11'b10110101010) ? 47'b00101011101110001011101010101111011101001000010 :
(key == 11'b10110101011) ? 47'b00101011101000101100111010101111010110101101101 :
(key == 11'b10110101100) ? 47'b00101011100011001110010010101111010000010011010 :
(key == 11'b10110101101) ? 47'b00101011011101101111111010101111001001111001011 :
(key == 11'b10110101110) ? 47'b00101011011000010001101010101111000011011111110 :
(key == 11'b10110101111) ? 47'b00101011010010110011101010101110111101000110100 :
(key == 11'b10110110000) ? 47'b00101011001101010101110010101110110110101101100 :
(key == 11'b10110110001) ? 47'b00101011000111111000001010101110110000010100111 :
(key == 11'b10110110010) ? 47'b00101011000010011010110010101110101001111100110 :
(key == 11'b10110110011) ? 47'b00101010111100111101101010101110100011100101000 :
(key == 11'b10110110100) ? 47'b00101010110111100000100010101110011101001101011 :
(key == 11'b10110110101) ? 47'b00101010110010000011110010101110010110110110010 :
(key == 11'b10110110110) ? 47'b00101010101100100111001010101110010000011111011 :
(key == 11'b10110110111) ? 47'b00101010100111001010110010101110001010001001000 :
(key == 11'b10110111000) ? 47'b00101010100001101110100010101110000011110010111 :
(key == 11'b10110111001) ? 47'b00101010011100010010100010101101111101011101001 :
(key == 11'b10110111010) ? 47'b00101010010110110110101010101101110111000111101 :
(key == 11'b10110111011) ? 47'b00101010010001011011000010101101110000110010100 :
(key == 11'b10110111100) ? 47'b00101010001011111111101010101101101010011101111 :
(key == 11'b10110111101) ? 47'b00101010000110100100011010101101100100001001011 :
(key == 11'b10110111110) ? 47'b00101010000001001001011010101101011101110101011 :
(key == 11'b10110111111) ? 47'b00101001111011101110100010101101010111100001101 :
(key == 11'b10111000000) ? 47'b00101001110110010011111010101101010001001110010 :
(key == 11'b10111000001) ? 47'b00101001110000111001011010101101001010111011010 :
(key == 11'b10111000010) ? 47'b00101001101011011111001010101101000100101000100 :
(key == 11'b10111000011) ? 47'b00101001100110000101001010101100111110010110010 :
(key == 11'b10111000100) ? 47'b00101001100000101011010010101100111000000100010 :
(key == 11'b10111000101) ? 47'b00101001011011010001101010101100110001110010101 :
(key == 11'b10111000110) ? 47'b00101001010101111000001010101100101011100001010 :
(key == 11'b10111000111) ? 47'b00101001010000011110111010101100100101010000011 :
(key == 11'b10111001000) ? 47'b00101001001011000101111010101100011110111111110 :
(key == 11'b10111001001) ? 47'b00101001000101101101000010101100011000101111100 :
(key == 11'b10111001010) ? 47'b00101001000000010100010010101100010010011111100 :
(key == 11'b10111001011) ? 47'b00101000111010111011111010101100001100010000000 :
(key == 11'b10111001100) ? 47'b00101000110101100011100010101100000110000000101 :
(key == 11'b10111001101) ? 47'b00101000110000001011100010101011111111110001110 :
(key == 11'b10111001110) ? 47'b00101000101010110011100010101011111001100011001 :
(key == 11'b10111001111) ? 47'b00101000100101011011111010101011110011010100111 :
(key == 11'b10111010000) ? 47'b00101000100000000100011010101011101101000111000 :
(key == 11'b10111010001) ? 47'b00101000011010101101000010101011100110111001011 :
(key == 11'b10111010010) ? 47'b00101000010101010101111010101011100000101100001 :
(key == 11'b10111010011) ? 47'b00101000001111111111000010101011011010011111010 :
(key == 11'b10111010100) ? 47'b00101000001010101000010010101011010100010010110 :
(key == 11'b10111010101) ? 47'b00101000000101010001110010101011001110000110100 :
(key == 11'b10111010110) ? 47'b00100111111111111011011010101011000111111010101 :
(key == 11'b10111010111) ? 47'b00100111111010100101010010101011000001101111001 :
(key == 11'b10111011000) ? 47'b00100111110101001111010010101010111011100011111 :
(key == 11'b10111011001) ? 47'b00100111101111111001100010101010110101011001000 :
(key == 11'b10111011010) ? 47'b00100111101010100011111010101010101111001110011 :
(key == 11'b10111011011) ? 47'b00100111100101001110100010101010101001000100001 :
(key == 11'b10111011100) ? 47'b00100111011111111001011010101010100010111010011 :
(key == 11'b10111011101) ? 47'b00100111011010100100011010101010011100110000110 :
(key == 11'b10111011110) ? 47'b00100111010101001111101010101010010110100111101 :
(key == 11'b10111011111) ? 47'b00100111001111111011000010101010010000011110110 :
(key == 11'b10111100000) ? 47'b00100111001010100110100010101010001010010110000 :
(key == 11'b10111100001) ? 47'b00100111000101010010010010101010000100001101110 :
(key == 11'b10111100010) ? 47'b00100110111111111110010010101001111110000110000 :
(key == 11'b10111100011) ? 47'b00100110111010101010011010101001110111111110011 :
(key == 11'b10111100100) ? 47'b00100110110101010110110010101001110001110111001 :
(key == 11'b10111100101) ? 47'b00100110110000000011010010101001101011110000010 :
(key == 11'b10111100110) ? 47'b00100110101010110000000010101001100101101001101 :
(key == 11'b10111100111) ? 47'b00100110100101011101000010101001011111100011100 :
(key == 11'b10111101000) ? 47'b00100110100000001010001010101001011001011101101 :
(key == 11'b10111101001) ? 47'b00100110011010110111011010101001010011011000000 :
(key == 11'b10111101010) ? 47'b00100110010101100100111010101001001101010010110 :
(key == 11'b10111101011) ? 47'b00100110010000010010100010101001000111001101110 :
(key == 11'b10111101100) ? 47'b00100110001011000000011010101001000001001001001 :
(key == 11'b10111101101) ? 47'b00100110000101101110100010101000111011000100111 :
(key == 11'b10111101110) ? 47'b00100110000000011100110010101000110101000001000 :
(key == 11'b10111101111) ? 47'b00100101111011001011001010101000101110111101010 :
(key == 11'b10111110000) ? 47'b00100101110101111001110010101000101000111010000 :
(key == 11'b10111110001) ? 47'b00100101110000101000101010101000100010110111001 :
(key == 11'b10111110010) ? 47'b00100101101011010111101010101000011100110100011 :
(key == 11'b10111110011) ? 47'b00100101100110000110110010101000010110110010000 :
(key == 11'b10111110100) ? 47'b00100101100000110110001010101000010000110000000 :
(key == 11'b10111110101) ? 47'b00100101011011100101110010101000001010101110011 :
(key == 11'b10111110110) ? 47'b00100101010110010101100010101000000100101101000 :
(key == 11'b10111110111) ? 47'b00100101010001000101100010100111111110101100001 :
(key == 11'b10111111000) ? 47'b00100101001011110101101010100111111000101011011 :
(key == 11'b10111111001) ? 47'b00100101000110100101111010100111110010101010111 :
(key == 11'b10111111010) ? 47'b00100101000001010110011010100111101100101010111 :
(key == 11'b10111111011) ? 47'b00100100111100000111001010100111100110101011001 :
(key == 11'b10111111100) ? 47'b00100100110110111000000010100111100000101011110 :
(key == 11'b10111111101) ? 47'b00100100110001101001001010100111011010101100110 :
(key == 11'b10111111110) ? 47'b00100100101100011010011010100111010100101101111 :
(key == 11'b10111111111) ? 47'b00100100100111001011110010100111001110101111011 :
(key == 11'b11000000000) ? 47'b00100100100001111101011010100111001000110001010 :
(key == 11'b11000000001) ? 47'b00100100011100101111010010100111000010110011100 :
(key == 11'b11000000010) ? 47'b00100100010111100001010010100110111100110110000 :
(key == 11'b11000000011) ? 47'b00100100010010010011011010100110110110111000110 :
(key == 11'b11000000100) ? 47'b00100100001101000101110010100110110000111011111 :
(key == 11'b11000000101) ? 47'b00100100000111111000011010100110101010111111011 :
(key == 11'b11000000110) ? 47'b00100100000010101011001010100110100101000011001 :
(key == 11'b11000000111) ? 47'b00100011111101011110000010100110011111000111010 :
(key == 11'b11000001000) ? 47'b00100011111000010001001010100110011001001011101 :
(key == 11'b11000001001) ? 47'b00100011110011000100100010100110010011010000011 :
(key == 11'b11000001010) ? 47'b00100011101101111000000010100110001101010101100 :
(key == 11'b11000001011) ? 47'b00100011101000101011101010100110000111011010110 :
(key == 11'b11000001100) ? 47'b00100011100011011111100010100110000001100000100 :
(key == 11'b11000001101) ? 47'b00100011011110010011100010100101111011100110011 :
(key == 11'b11000001110) ? 47'b00100011011001000111110010100101110101101100110 :
(key == 11'b11000001111) ? 47'b00100011010011111100010010100101101111110011100 :
(key == 11'b11000010000) ? 47'b00100011001110110000110010100101101001111010010 :
(key == 11'b11000010001) ? 47'b00100011001001100101101010100101100100000001101 :
(key == 11'b11000010010) ? 47'b00100011000100011010100010100101011110001001001 :
(key == 11'b11000010011) ? 47'b00100010111111001111110010100101011000010001001 :
(key == 11'b11000010100) ? 47'b00100010111010000101000010100101010010011001010 :
(key == 11'b11000010101) ? 47'b00100010110100111010100010100101001100100001110 :
(key == 11'b11000010110) ? 47'b00100010101111110000010010100101000110101010101 :
(key == 11'b11000010111) ? 47'b00100010101010100110001010100101000000110011110 :
(key == 11'b11000011000) ? 47'b00100010100101011100010010100100111010111101010 :
(key == 11'b11000011001) ? 47'b00100010100000010010100010100100110101000111000 :
(key == 11'b11000011010) ? 47'b00100010011011001000111010100100101111010001000 :
(key == 11'b11000011011) ? 47'b00100010010101111111100010100100101001011011011 :
(key == 11'b11000011100) ? 47'b00100010010000110110010010100100100011100110000 :
(key == 11'b11000011101) ? 47'b00100010001011101101010010100100011101110001000 :
(key == 11'b11000011110) ? 47'b00100010000110100100011010100100010111111100010 :
(key == 11'b11000011111) ? 47'b00100010000001011011110010100100010010000111111 :
(key == 11'b11000100000) ? 47'b00100001111100010011010010100100001100010011110 :
(key == 11'b11000100001) ? 47'b00100001110111001011000010100100000110100000001 :
(key == 11'b11000100010) ? 47'b00100001110010000010111010100100000000101100101 :
(key == 11'b11000100011) ? 47'b00100001101100111011000010100011111010111001100 :
(key == 11'b11000100100) ? 47'b00100001100111110011010010100011110101000110101 :
(key == 11'b11000100101) ? 47'b00100001100010101011101010100011101111010100001 :
(key == 11'b11000100110) ? 47'b00100001011101100100010010100011101001100001111 :
(key == 11'b11000100111) ? 47'b00100001011000011101000010100011100011101111111 :
(key == 11'b11000101000) ? 47'b00100001010011010110000010100011011101111110010 :
(key == 11'b11000101001) ? 47'b00100001001110001111001010100011011000001101000 :
(key == 11'b11000101010) ? 47'b00100001001001001000100010100011010010011100000 :
(key == 11'b11000101011) ? 47'b00100001000100000010000010100011001100101011010 :
(key == 11'b11000101100) ? 47'b00100000111110111011110010100011000110111010111 :
(key == 11'b11000101101) ? 47'b00100000111001110101101010100011000001001010111 :
(key == 11'b11000101110) ? 47'b00100000110100101111101010100010111011011011000 :
(key == 11'b11000101111) ? 47'b00100000101111101001111010100010110101101011100 :
(key == 11'b11000110000) ? 47'b00100000101010100100010010100010101111111100010 :
(key == 11'b11000110001) ? 47'b00100000100101011110111010100010101010001101100 :
(key == 11'b11000110010) ? 47'b00100000100000011001101010100010100100011110111 :
(key == 11'b11000110011) ? 47'b00100000011011010100101010100010011110110000101 :
(key == 11'b11000110100) ? 47'b00100000010110001111110010100010011001000010101 :
(key == 11'b11000110101) ? 47'b00100000010001001011000010100010010011010100111 :
(key == 11'b11000110110) ? 47'b00100000001100000110100010100010001101100111101 :
(key == 11'b11000110111) ? 47'b00100000000111000010001010100010000111111010100 :
(key == 11'b11000111000) ? 47'b00100000000001111110000010100010000010001101110 :
(key == 11'b11000111001) ? 47'b00011111111100111010000010100001111100100001010 :
(key == 11'b11000111010) ? 47'b00011111110111110110010010100001110110110101001 :
(key == 11'b11000111011) ? 47'b00011111110010110010101010100001110001001001010 :
(key == 11'b11000111100) ? 47'b00011111101101101111001010100001101011011101101 :
(key == 11'b11000111101) ? 47'b00011111101000101011111010100001100101110010011 :
(key == 11'b11000111110) ? 47'b00011111100011101000110010100001100000000111011 :
(key == 11'b11000111111) ? 47'b00011111011110100101111010100001011010011100110 :
(key == 11'b11001000000) ? 47'b00011111011001100011001010100001010100110010011 :
(key == 11'b11001000001) ? 47'b00011111010100100000101010100001001111001000011 :
(key == 11'b11001000010) ? 47'b00011111001111011110010010100001001001011110101 :
(key == 11'b11001000011) ? 47'b00011111001010011100000010100001000011110101001 :
(key == 11'b11001000100) ? 47'b00011111000101011010000010100000111110001011111 :
(key == 11'b11001000101) ? 47'b00011111000000011000001010100000111000100011000 :
(key == 11'b11001000110) ? 47'b00011110111011010110011010100000110010111010011 :
(key == 11'b11001000111) ? 47'b00011110110110010100111010100000101101010010000 :
(key == 11'b11001001000) ? 47'b00011110110001010011101010100000100111101010001 :
(key == 11'b11001001001) ? 47'b00011110101100010010100010100000100010000010100 :
(key == 11'b11001001010) ? 47'b00011110100111010001100010100000011100011011000 :
(key == 11'b11001001011) ? 47'b00011110100010010000101010100000010110110011111 :
(key == 11'b11001001100) ? 47'b00011110011101010000000010100000010001001101000 :
(key == 11'b11001001101) ? 47'b00011110011000001111101010100000001011100110101 :
(key == 11'b11001001110) ? 47'b00011110010011001111011010100000000110000000011 :
(key == 11'b11001001111) ? 47'b00011110001110001111010010100000000000011010011 :
(key == 11'b11001010000) ? 47'b00011110001001001111010010011111111010110100101 :
(key == 11'b11001010001) ? 47'b00011110000100001111100010011111110101001111011 :
(key == 11'b11001010010) ? 47'b00011101111111010000000010011111101111101010011 :
(key == 11'b11001010011) ? 47'b00011101111010010000100010011111101010000101100 :
(key == 11'b11001010100) ? 47'b00011101110101010001011010011111100100100001001 :
(key == 11'b11001010101) ? 47'b00011101110000010010010010011111011110111100111 :
(key == 11'b11001010110) ? 47'b00011101101011010011011010011111011001011001000 :
(key == 11'b11001010111) ? 47'b00011101100110010100110010011111010011110101100 :
(key == 11'b11001011000) ? 47'b00011101100001010110001010011111001110010010000 :
(key == 11'b11001011001) ? 47'b00011101011100010111110010011111001000101111000 :
(key == 11'b11001011010) ? 47'b00011101010111011001101010011111000011001100011 :
(key == 11'b11001011011) ? 47'b00011101010010011011101010011110111101101001111 :
(key == 11'b11001011100) ? 47'b00011101001101011101110010011110111000000111110 :
(key == 11'b11001011101) ? 47'b00011101001000100000001010011110110010100101111 :
(key == 11'b11001011110) ? 47'b00011101000011100010101010011110101101000100010 :
(key == 11'b11001011111) ? 47'b00011100111110100101010010011110100111100011000 :
(key == 11'b11001100000) ? 47'b00011100111001101000001010011110100010000010000 :
(key == 11'b11001100001) ? 47'b00011100110100101011001010011110011100100001010 :
(key == 11'b11001100010) ? 47'b00011100101111101110011010011110010111000000111 :
(key == 11'b11001100011) ? 47'b00011100101010110001110010011110010001100000110 :
(key == 11'b11001100100) ? 47'b00011100100101110101010010011110001100000000111 :
(key == 11'b11001100101) ? 47'b00011100100000111001000010011110000110100001011 :
(key == 11'b11001100110) ? 47'b00011100011011111100111010011110000001000010000 :
(key == 11'b11001100111) ? 47'b00011100010111000000111010011101111011100011000 :
(key == 11'b11001101000) ? 47'b00011100010010000101001010011101110110000100010 :
(key == 11'b11001101001) ? 47'b00011100001101001001100010011101110000100101111 :
(key == 11'b11001101010) ? 47'b00011100001000001110001010011101101011000111110 :
(key == 11'b11001101011) ? 47'b00011100000011010010111010011101100101101001111 :
(key == 11'b11001101100) ? 47'b00011011111110010111110010011101100000001100011 :
(key == 11'b11001101101) ? 47'b00011011111001011100110010011101011010101111000 :
(key == 11'b11001101110) ? 47'b00011011110100100010000010011101010101010010000 :
(key == 11'b11001101111) ? 47'b00011011101111100111100010011101001111110101011 :
(key == 11'b11001110000) ? 47'b00011011101010101101001010011101001010011000111 :
(key == 11'b11001110001) ? 47'b00011011100101110010111010011101000100111100110 :
(key == 11'b11001110010) ? 47'b00011011100000111000110010011100111111100000111 :
(key == 11'b11001110011) ? 47'b00011011011011111110111010011100111010000101010 :
(key == 11'b11001110100) ? 47'b00011011010111000101001010011100110100101001111 :
(key == 11'b11001110101) ? 47'b00011011010010001011101010011100101111001111000 :
(key == 11'b11001110110) ? 47'b00011011001101010010001010011100101001110100001 :
(key == 11'b11001110111) ? 47'b00011011001000011001000010011100100100011001110 :
(key == 11'b11001111000) ? 47'b00011011000011011111111010011100011110111111100 :
(key == 11'b11001111001) ? 47'b00011010111110100111000010011100011001100101101 :
(key == 11'b11001111010) ? 47'b00011010111001101110010010011100010100001011111 :
(key == 11'b11001111011) ? 47'b00011010110100110101110010011100001110110010101 :
(key == 11'b11001111100) ? 47'b00011010101111111101011010011100001001011001101 :
(key == 11'b11001111101) ? 47'b00011010101011000101001010011100000100000000110 :
(key == 11'b11001111110) ? 47'b00011010100110001101001010011011111110101000010 :
(key == 11'b11001111111) ? 47'b00011010100001010101010010011011111001010000000 :
(key == 11'b11010000000) ? 47'b00011010011100011101100010011011110011111000000 :
(key == 11'b11010000001) ? 47'b00011010010111100110000010011011101110100000011 :
(key == 11'b11010000010) ? 47'b00011010010010101110101010011011101001001001000 :
(key == 11'b11010000011) ? 47'b00011010001101110111100010011011100011110010000 :
(key == 11'b11010000100) ? 47'b00011010001001000000011010011011011110011011000 :
(key == 11'b11010000101) ? 47'b00011010000100001001100010011011011001000100100 :
(key == 11'b11010000110) ? 47'b00011001111111010010111010011011010011101110010 :
(key == 11'b11010000111) ? 47'b00011001111010011100010010011011001110011000001 :
(key == 11'b11010001000) ? 47'b00011001110101100110000010011011001001000010100 :
(key == 11'b11010001001) ? 47'b00011001110000101111110010011011000011101101000 :
(key == 11'b11010001010) ? 47'b00011001101011111001110010011010111110010111111 :
(key == 11'b11010001011) ? 47'b00011001100111000011111010011010111001000011000 :
(key == 11'b11010001100) ? 47'b00011001100010001110001010011010110011101110010 :
(key == 11'b11010001101) ? 47'b00011001011101011000101010011010101110011001111 :
(key == 11'b11010001110) ? 47'b00011001011000100011010010011010101001000101111 :
(key == 11'b11010001111) ? 47'b00011001010011101110000010011010100011110010000 :
(key == 11'b11010010000) ? 47'b00011001001110111001000010011010011110011110100 :
(key == 11'b11010010001) ? 47'b00011001001010000100001010011010011001001011010 :
(key == 11'b11010010010) ? 47'b00011001000101001111011010011010010011111000001 :
(key == 11'b11010010011) ? 47'b00011001000000011010111010011010001110100101100 :
(key == 11'b11010010100) ? 47'b00011000111011100110100010011010001001010011000 :
(key == 11'b11010010101) ? 47'b00011000110110110010010010011010000100000000110 :
(key == 11'b11010010110) ? 47'b00011000110001111110010010011001111110101110111 :
(key == 11'b11010010111) ? 47'b00011000101101001010011010011001111001011101010 :
(key == 11'b11010011000) ? 47'b00011000101000010110101010011001110100001011111 :
(key == 11'b11010011001) ? 47'b00011000100011100011001010011001101110111010111 :
(key == 11'b11010011010) ? 47'b00011000011110101111110010011001101001101010000 :
(key == 11'b11010011011) ? 47'b00011000011001111100100010011001100100011001100 :
(key == 11'b11010011100) ? 47'b00011000010101001001100010011001011111001001010 :
(key == 11'b11010011101) ? 47'b00011000010000010110101010011001011001111001010 :
(key == 11'b11010011110) ? 47'b00011000001011100011111010011001010100101001100 :
(key == 11'b11010011111) ? 47'b00011000000110110001010010011001001111011001111 :
(key == 11'b11010100000) ? 47'b00011000000001111110111010011001001010001010110 :
(key == 11'b11010100001) ? 47'b00010111111101001100101010011001000100111011110 :
(key == 11'b11010100010) ? 47'b00010111111000011010101010011000111111101101010 :
(key == 11'b11010100011) ? 47'b00010111110011101000101010011000111010011110110 :
(key == 11'b11010100100) ? 47'b00010111101110110110111010011000110101010000100 :
(key == 11'b11010100101) ? 47'b00010111101010000101011010011000110000000010110 :
(key == 11'b11010100110) ? 47'b00010111100101010011111010011000101010110101001 :
(key == 11'b11010100111) ? 47'b00010111100000100010101010011000100101100111110 :
(key == 11'b11010101000) ? 47'b00010111011011110001101010011000100000011010110 :
(key == 11'b11010101001) ? 47'b00010111010111000000101010011000011011001101111 :
(key == 11'b11010101010) ? 47'b00010111010010001111111010011000010110000001011 :
(key == 11'b11010101011) ? 47'b00010111001101011111010010011000010000110101001 :
(key == 11'b11010101100) ? 47'b00010111001000101110111010011000001011101001010 :
(key == 11'b11010101101) ? 47'b00010111000011111110100010011000000110011101011 :
(key == 11'b11010101110) ? 47'b00010110111111001110011010011000000001010001111 :
(key == 11'b11010101111) ? 47'b00010110111010011110100010010111111100000110110 :
(key == 11'b11010110000) ? 47'b00010110110101101110101010010111110110111011110 :
(key == 11'b11010110001) ? 47'b00010110110000111111000010010111110001110001001 :
(key == 11'b11010110010) ? 47'b00010110101100001111100010010111101100100110101 :
(key == 11'b11010110011) ? 47'b00010110100111100000010010010111100111011100100 :
(key == 11'b11010110100) ? 47'b00010110100010110001001010010111100010010010101 :
(key == 11'b11010110101) ? 47'b00010110011110000010001010010111011101001001000 :
(key == 11'b11010110110) ? 47'b00010110011001010011010010010111010111111111101 :
(key == 11'b11010110111) ? 47'b00010110010100100100101010010111010010110110101 :
(key == 11'b11010111000) ? 47'b00010110001111110110001010010111001101101101110 :
(key == 11'b11010111001) ? 47'b00010110001011000111110010010111001000100101001 :
(key == 11'b11010111010) ? 47'b00010110000110011001100010010111000011011100110 :
(key == 11'b11010111011) ? 47'b00010110000001101011100010010110111110010100110 :
(key == 11'b11010111100) ? 47'b00010101111100111101101010010110111001001100111 :
(key == 11'b11010111101) ? 47'b00010101111000010000000010010110110100000101100 :
(key == 11'b11010111110) ? 47'b00010101110011100010011010010110101110111110001 :
(key == 11'b11010111111) ? 47'b00010101101110110101000010010110101001110111001 :
(key == 11'b11011000000) ? 47'b00010101101010000111110010010110100100110000011 :
(key == 11'b11011000001) ? 47'b00010101100101011010110010010110011111101001111 :
(key == 11'b11011000010) ? 47'b00010101100000101101110010010110011010100011100 :
(key == 11'b11011000011) ? 47'b00010101011100000001000010010110010101011101101 :
(key == 11'b11011000100) ? 47'b00010101010111010100100010010110010000011000000 :
(key == 11'b11011000101) ? 47'b00010101010010101000000010010110001011010010011 :
(key == 11'b11011000110) ? 47'b00010101001101111011110010010110000110001101010 :
(key == 11'b11011000111) ? 47'b00010101001001001111101010010110000001001000010 :
(key == 11'b11011001000) ? 47'b00010101000100100011101010010101111100000011100 :
(key == 11'b11011001001) ? 47'b00010100111111110111111010010101110110111111001 :
(key == 11'b11011001010) ? 47'b00010100111011001100010010010101110001111011000 :
(key == 11'b11011001011) ? 47'b00010100110110100000110010010101101100110111001 :
(key == 11'b11011001100) ? 47'b00010100110001110101100010010101100111110011100 :
(key == 11'b11011001101) ? 47'b00010100101101001010010010010101100010110000000 :
(key == 11'b11011001110) ? 47'b00010100101000011111010010010101011101101100111 :
(key == 11'b11011001111) ? 47'b00010100100011110100011010010101011000101010000 :
(key == 11'b11011010000) ? 47'b00010100011111001001110010010101010011100111011 :
(key == 11'b11011010001) ? 47'b00010100011010011111010010010101001110100101000 :
(key == 11'b11011010010) ? 47'b00010100010101110100111010010101001001100010111 :
(key == 11'b11011010011) ? 47'b00010100010001001010101010010101000100100001000 :
(key == 11'b11011010100) ? 47'b00010100001100100000100010010100111111011111011 :
(key == 11'b11011010101) ? 47'b00010100000111110110101010010100111010011110000 :
(key == 11'b11011010110) ? 47'b00010100000011001100111010010100110101011100111 :
(key == 11'b11011010111) ? 47'b00010011111110100011010010010100110000011100000 :
(key == 11'b11011011000) ? 47'b00010011111001111001111010010100101011011011100 :
(key == 11'b11011011001) ? 47'b00010011110101010000101010010100100110011011001 :
(key == 11'b11011011010) ? 47'b00010011110000100111100010010100100001011011000 :
(key == 11'b11011011011) ? 47'b00010011101011111110100010010100011100011011001 :
(key == 11'b11011011100) ? 47'b00010011100111010101101010010100010111011011100 :
(key == 11'b11011011101) ? 47'b00010011100010101101000010010100010010011100001 :
(key == 11'b11011011110) ? 47'b00010011011110000100100010010100001101011101001 :
(key == 11'b11011011111) ? 47'b00010011011001011100001010010100001000011110010 :
(key == 11'b11011100000) ? 47'b00010011010100110100000010010100000011011111101 :
(key == 11'b11011100001) ? 47'b00010011010000001100000010010011111110100001011 :
(key == 11'b11011100010) ? 47'b00010011001011100100001010010011111001100011010 :
(key == 11'b11011100011) ? 47'b00010011000110111100011010010011110100100101011 :
(key == 11'b11011100100) ? 47'b00010011000010010100110010010011101111100111110 :
(key == 11'b11011100101) ? 47'b00010010111101101101011010010011101010101010100 :
(key == 11'b11011100110) ? 47'b00010010111001000110001010010011100101101101011 :
(key == 11'b11011100111) ? 47'b00010010110100011111000010010011100000110000100 :
(key == 11'b11011101000) ? 47'b00010010101111111000001010010011011011110100000 :
(key == 11'b11011101001) ? 47'b00010010101011010001010010010011010110110111101 :
(key == 11'b11011101010) ? 47'b00010010100110101010101010010011010001111011100 :
(key == 11'b11011101011) ? 47'b00010010100010000100001010010011001100111111101 :
(key == 11'b11011101100) ? 47'b00010010011101011101111010010011001000000100001 :
(key == 11'b11011101101) ? 47'b00010010011000110111101010010011000011001000110 :
(key == 11'b11011101110) ? 47'b00010010010100010001101010010010111110001101101 :
(key == 11'b11011101111) ? 47'b00010010001111101011110010010010111001010010110 :
(key == 11'b11011110000) ? 47'b00010010001011000110001010010010110100011000010 :
(key == 11'b11011110001) ? 47'b00010010000110100000100010010010101111011101111 :
(key == 11'b11011110010) ? 47'b00010010000001111011001010010010101010100011110 :
(key == 11'b11011110011) ? 47'b00010001111101010101111010010010100101101001111 :
(key == 11'b11011110100) ? 47'b00010001111000110000110010010010100000110000010 :
(key == 11'b11011110101) ? 47'b00010001110100001011110010010010011011110110111 :
(key == 11'b11011110110) ? 47'b00010001101111100111000010010010010110111101110 :
(key == 11'b11011110111) ? 47'b00010001101011000010011010010010010010000100111 :
(key == 11'b11011111000) ? 47'b00010001100110011101111010010010001101001100010 :
(key == 11'b11011111001) ? 47'b00010001100001111001100010010010001000010011110 :
(key == 11'b11011111010) ? 47'b00010001011101010101011010010010000011011011110 :
(key == 11'b11011111011) ? 47'b00010001011000110001011010010001111110100011111 :
(key == 11'b11011111100) ? 47'b00010001010100001101100010010001111001101100001 :
(key == 11'b11011111101) ? 47'b00010001001111101001110010010001110100110100110 :
(key == 11'b11011111110) ? 47'b00010001001011000110001010010001101111111101100 :
(key == 11'b11011111111) ? 47'b00010001000110100010110010010001101011000110101 :
(key == 11'b11100000000) ? 47'b00010001000001111111100010010001100110010000000 :
(key == 11'b11100000001) ? 47'b00010000111101011100011010010001100001011001100 :
(key == 11'b11100000010) ? 47'b00010000111000111001011010010001011100100011010 :
(key == 11'b11100000011) ? 47'b00010000110100010110100010010001010111101101010 :
(key == 11'b11100000100) ? 47'b00010000101111110011111010010001010010110111100 :
(key == 11'b11100000101) ? 47'b00010000101011010001011010010001001110000010001 :
(key == 11'b11100000110) ? 47'b00010000100110101111000010010001001001001100111 :
(key == 11'b11100000111) ? 47'b00010000100010001100110010010001000100010111110 :
(key == 11'b11100001000) ? 47'b00010000011101101010110010010000111111100011001 :
(key == 11'b11100001001) ? 47'b00010000011001001000111010010000111010101110101 :
(key == 11'b11100001010) ? 47'b00010000010100100111000010010000110101111010010 :
(key == 11'b11100001011) ? 47'b00010000010000000101100010010000110001000110011 :
(key == 11'b11100001100) ? 47'b00010000001011100100000010010000101100010010100 :
(key == 11'b11100001101) ? 47'b00010000000111000010101010010000100111011110111 :
(key == 11'b11100001110) ? 47'b00010000000010100001100010010000100010101011101 :
(key == 11'b11100001111) ? 47'b00001111111110000000100010010000011101111000100 :
(key == 11'b11100010000) ? 47'b00001111111001011111101010010000011001000101101 :
(key == 11'b11100010001) ? 47'b00001111110100111111000010010000010100010011001 :
(key == 11'b11100010010) ? 47'b00001111110000011110011010010000001111100000110 :
(key == 11'b11100010011) ? 47'b00001111101011111110000010010000001010101110101 :
(key == 11'b11100010100) ? 47'b00001111100111011101110010010000000101111100110 :
(key == 11'b11100010101) ? 47'b00001111100010111101101010010000000001001011001 :
(key == 11'b11100010110) ? 47'b00001111011110011101101010001111111100011001101 :
(key == 11'b11100010111) ? 47'b00001111011001111101111010001111110111101000100 :
(key == 11'b11100011000) ? 47'b00001111010101011110001010001111110010110111100 :
(key == 11'b11100011001) ? 47'b00001111010000111110101010001111101110000110111 :
(key == 11'b11100011010) ? 47'b00001111001100011111010010001111101001010110011 :
(key == 11'b11100011011) ? 47'b00001111001000000000001010001111100100100110010 :
(key == 11'b11100011100) ? 47'b00001111000011100001000010001111011111110110001 :
(key == 11'b11100011101) ? 47'b00001110111111000010001010001111011011000110100 :
(key == 11'b11100011110) ? 47'b00001110111010100011010010001111010110010110111 :
(key == 11'b11100011111) ? 47'b00001110110110000100101010001111010001100111100 :
(key == 11'b11100100000) ? 47'b00001110110001100110010010001111001100111000101 :
(key == 11'b11100100001) ? 47'b00001110101101000111111010001111001000001001110 :
(key == 11'b11100100010) ? 47'b00001110101000101001110010001111000011011011010 :
(key == 11'b11100100011) ? 47'b00001110100100001011101010001110111110101100110 :
(key == 11'b11100100100) ? 47'b00001110011111101101110010001110111001111110101 :
(key == 11'b11100100101) ? 47'b00001110011011010000000010001110110101010000110 :
(key == 11'b11100100110) ? 47'b00001110010110110010100010001110110000100011010 :
(key == 11'b11100100111) ? 47'b00001110010010010101000010001110101011110101110 :
(key == 11'b11100101000) ? 47'b00001110001101110111110010001110100111001000101 :
(key == 11'b11100101001) ? 47'b00001110001001011010100010001110100010011011101 :
(key == 11'b11100101010) ? 47'b00001110000100111101100010001110011101101110111 :
(key == 11'b11100101011) ? 47'b00001110000000100000110010001110011001000010100 :
(key == 11'b11100101100) ? 47'b00001101111100000100000010001110010100010110010 :
(key == 11'b11100101101) ? 47'b00001101110111100111011010001110001111101010001 :
(key == 11'b11100101110) ? 47'b00001101110011001011000010001110001010111110011 :
(key == 11'b11100101111) ? 47'b00001101101110101110110010001110000110010010111 :
(key == 11'b11100110000) ? 47'b00001101101010010010101010001110000001100111100 :
(key == 11'b11100110001) ? 47'b00001101100101110110101010001101111100111100011 :
(key == 11'b11100110010) ? 47'b00001101100001011010110010001101111000010001100 :
(key == 11'b11100110011) ? 47'b00001101011100111111001010001101110011100111000 :
(key == 11'b11100110100) ? 47'b00001101011000100011101010001101101110111100101 :
(key == 11'b11100110101) ? 47'b00001101010100001000001010001101101010010010010 :
(key == 11'b11100110110) ? 47'b00001101001111101100111010001101100101101000011 :
(key == 11'b11100110111) ? 47'b00001101001011010001111010001101100000111110110 :
(key == 11'b11100111000) ? 47'b00001101000110110110111010001101011100010101010 :
(key == 11'b11100111001) ? 47'b00001101000010011100001010001101010111101100000 :
(key == 11'b11100111010) ? 47'b00001100111110000001011010001101010011000010111 :
(key == 11'b11100111011) ? 47'b00001100111001100110111010001101001110011010001 :
(key == 11'b11100111100) ? 47'b00001100110101001100100010001101001001110001101 :
(key == 11'b11100111101) ? 47'b00001100110000110010010010001101000101001001010 :
(key == 11'b11100111110) ? 47'b00001100101100011000001010001101000000100001001 :
(key == 11'b11100111111) ? 47'b00001100100111111110010010001100111011111001010 :
(key == 11'b11101000000) ? 47'b00001100100011100100011010001100110111010001100 :
(key == 11'b11101000001) ? 47'b00001100011111001010110010001100110010101010001 :
(key == 11'b11101000010) ? 47'b00001100011010110001010010001100101110000010111 :
(key == 11'b11101000011) ? 47'b00001100010110010111111010001100101001011100000 :
(key == 11'b11101000100) ? 47'b00001100010001111110101010001100100100110101001 :
(key == 11'b11101000101) ? 47'b00001100001101100101101010001100100000001110110 :
(key == 11'b11101000110) ? 47'b00001100001001001100101010001100011011101000011 :
(key == 11'b11101000111) ? 47'b00001100000100110011111010001100010111000010011 :
(key == 11'b11101001000) ? 47'b00001100000000011011010010001100010010011100100 :
(key == 11'b11101001001) ? 47'b00001011111100000010110010001100001101110110111 :
(key == 11'b11101001010) ? 47'b00001011110111101010011010001100001001010001100 :
(key == 11'b11101001011) ? 47'b00001011110011010010001010001100000100101100010 :
(key == 11'b11101001100) ? 47'b00001011101110111010000010001100000000000111010 :
(key == 11'b11101001101) ? 47'b00001011101010100010001010001011111011100010101 :
(key == 11'b11101001110) ? 47'b00001011100110001010011010001011110110111110001 :
(key == 11'b11101001111) ? 47'b00001011100001110010110010001011110010011001111 :
(key == 11'b11101010000) ? 47'b00001011011101011011010010001011101101110101111 :
(key == 11'b11101010001) ? 47'b00001011011001000011111010001011101001010010000 :
(key == 11'b11101010010) ? 47'b00001011010100101100101010001011100100101110011 :
(key == 11'b11101010011) ? 47'b00001011010000010101100010001011100000001010111 :
(key == 11'b11101010100) ? 47'b00001011001011111110101010001011011011100111111 :
(key == 11'b11101010101) ? 47'b00001011000111100111110010001011010111000100110 :
(key == 11'b11101010110) ? 47'b00001011000011010001001010001011010010100010001 :
(key == 11'b11101010111) ? 47'b00001010111110111010101010001011001101111111101 :
(key == 11'b11101011000) ? 47'b00001010111010100100010010001011001001011101011 :
(key == 11'b11101011001) ? 47'b00001010110110001110000010001011000100111011010 :
(key == 11'b11101011010) ? 47'b00001010110001111000000010001011000000011001100 :
(key == 11'b11101011011) ? 47'b00001010101101100010000010001010111011110111111 :
(key == 11'b11101011100) ? 47'b00001010101001001100010010001010110111010110100 :
(key == 11'b11101011101) ? 47'b00001010100100110110101010001010110010110101011 :
(key == 11'b11101011110) ? 47'b00001010100000100001000010001010101110010100011 :
(key == 11'b11101011111) ? 47'b00001010011100001011101010001010101001110011101 :
(key == 11'b11101100000) ? 47'b00001010010111110110100010001010100101010011010 :
(key == 11'b11101100001) ? 47'b00001010010011100001011010001010100000110010111 :
(key == 11'b11101100010) ? 47'b00001010001111001100011010001010011100010010110 :
(key == 11'b11101100011) ? 47'b00001010001010110111101010001010010111110011000 :
(key == 11'b11101100100) ? 47'b00001010000110100010111010001010010011010011010 :
(key == 11'b11101100101) ? 47'b00001010000010001110011010001010001110110011111 :
(key == 11'b11101100110) ? 47'b00001001111101111010000010001010001010010100110 :
(key == 11'b11101100111) ? 47'b00001001111001100101110010001010000101110101110 :
(key == 11'b11101101000) ? 47'b00001001110101010001101010001010000001010111000 :
(key == 11'b11101101001) ? 47'b00001001110000111101101010001001111100111000100 :
(key == 11'b11101101010) ? 47'b00001001101100101001110010001001111000011010001 :
(key == 11'b11101101011) ? 47'b00001001101000010110001010001001110011111100000 :
(key == 11'b11101101100) ? 47'b00001001100100000010100010001001101111011110001 :
(key == 11'b11101101101) ? 47'b00001001011111101111001010001001101011000000100 :
(key == 11'b11101101110) ? 47'b00001001011011011011111010001001100110100011000 :
(key == 11'b11101101111) ? 47'b00001001010111001000110010001001100010000101111 :
(key == 11'b11101110000) ? 47'b00001001010010110101110010001001011101101000110 :
(key == 11'b11101110001) ? 47'b00001001001110100010111010001001011001001100000 :
(key == 11'b11101110010) ? 47'b00001001001010010000001010001001010100101111011 :
(key == 11'b11101110011) ? 47'b00001001000101111101101010001001010000010011001 :
(key == 11'b11101110100) ? 47'b00001001000001101011001010001001001011110110111 :
(key == 11'b11101110101) ? 47'b00001000111101011000111010001001000111011011000 :
(key == 11'b11101110110) ? 47'b00001000111001000110101010001001000010111111001 :
(key == 11'b11101110111) ? 47'b00001000110100110100101010001000111110100011110 :
(key == 11'b11101111000) ? 47'b00001000110000100010110010001000111010001000011 :
(key == 11'b11101111001) ? 47'b00001000101100010001000010001000110101101101011 :
(key == 11'b11101111010) ? 47'b00001000100111111111011010001000110001010010100 :
(key == 11'b11101111011) ? 47'b00001000100011101110000010001000101100110111111 :
(key == 11'b11101111100) ? 47'b00001000011111011100101010001000101000011101011 :
(key == 11'b11101111101) ? 47'b00001000011011001011011010001000100100000011001 :
(key == 11'b11101111110) ? 47'b00001000010110111010011010001000011111101001010 :
(key == 11'b11101111111) ? 47'b00001000010010101001100010001000011011001111100 :
(key == 11'b11110000000) ? 47'b00001000001110011000101010001000010110110101110 :
(key == 11'b11110000001) ? 47'b00001000001010001000000010001000010010011100011 :
(key == 11'b11110000010) ? 47'b00001000000101110111100010001000001110000011010 :
(key == 11'b11110000011) ? 47'b00001000000001100111001010001000001001101010011 :
(key == 11'b11110000100) ? 47'b00000111111101010110111010001000000101010001101 :
(key == 11'b11110000101) ? 47'b00000111111001000110110010001000000000111001000 :
(key == 11'b11110000110) ? 47'b00000111110100110110111010000111111100100000110 :
(key == 11'b11110000111) ? 47'b00000111110000100111000010000111111000001000101 :
(key == 11'b11110001000) ? 47'b00000111101100010111011010000111110011110000111 :
(key == 11'b11110001001) ? 47'b00000111101000000111110010000111101111011001001 :
(key == 11'b11110001010) ? 47'b00000111100011111000011010000111101011000001101 :
(key == 11'b11110001011) ? 47'b00000111011111101001001010000111100110101010011 :
(key == 11'b11110001100) ? 47'b00000111011011011010000010000111100010010011011 :
(key == 11'b11110001101) ? 47'b00000111010111001011000010000111011101111100101 :
(key == 11'b11110001110) ? 47'b00000111010010111100001010000111011001100110000 :
(key == 11'b11110001111) ? 47'b00000111001110101101011010000111010101001111100 :
(key == 11'b11110010000) ? 47'b00000111001010011110110010000111010000111001010 :
(key == 11'b11110010001) ? 47'b00000111000110010000010010000111001100100011010 :
(key == 11'b11110010010) ? 47'b00000111000010000010000010000111001000001101100 :
(key == 11'b11110010011) ? 47'b00000110111101110011110010000111000011110111111 :
(key == 11'b11110010100) ? 47'b00000110111001100101110010000110111111100010101 :
(key == 11'b11110010101) ? 47'b00000110110101010111111010000110111011001101100 :
(key == 11'b11110010110) ? 47'b00000110110001001010000010000110110110111000011 :
(key == 11'b11110010111) ? 47'b00000110101100111100011010000110110010100011110 :
(key == 11'b11110011000) ? 47'b00000110101000101110111010000110101110001111001 :
(key == 11'b11110011001) ? 47'b00000110100100100001100010000110101001111010111 :
(key == 11'b11110011010) ? 47'b00000110100000010100010010000110100101100110110 :
(key == 11'b11110011011) ? 47'b00000110011100000111001010000110100001010010110 :
(key == 11'b11110011100) ? 47'b00000110010111111010001010000110011100111111001 :
(key == 11'b11110011101) ? 47'b00000110010011101101011010000110011000101011101 :
(key == 11'b11110011110) ? 47'b00000110001111100000101010000110010100011000011 :
(key == 11'b11110011111) ? 47'b00000110001011010100000010000110010000000101001 :
(key == 11'b11110100000) ? 47'b00000110000111000111101010000110001011110010011 :
(key == 11'b11110100001) ? 47'b00000110000010111011011010000110000111011111110 :
(key == 11'b11110100010) ? 47'b00000101111110101111001010000110000011001101010 :
(key == 11'b11110100011) ? 47'b00000101111010100011001010000101111110111011000 :
(key == 11'b11110100100) ? 47'b00000101110110010111010010000101111010101001000 :
(key == 11'b11110100101) ? 47'b00000101110010001011100010000101110110010111001 :
(key == 11'b11110100110) ? 47'b00000101101101111111111010000101110010000101100 :
(key == 11'b11110100111) ? 47'b00000101101001110100011010000101101101110100000 :
(key == 11'b11110101000) ? 47'b00000101100101101001000010000101101001100010110 :
(key == 11'b11110101001) ? 47'b00000101100001011101110010000101100101010001110 :
(key == 11'b11110101010) ? 47'b00000101011101010010101010000101100001000000111 :
(key == 11'b11110101011) ? 47'b00000101011001000111101010000101011100110000010 :
(key == 11'b11110101100) ? 47'b00000101010100111100111010000101011000011111111 :
(key == 11'b11110101101) ? 47'b00000101010000110010001010000101010100001111101 :
(key == 11'b11110101110) ? 47'b00000101001100100111101010000101001111111111101 :
(key == 11'b11110101111) ? 47'b00000101001000011101001010000101001011101111110 :
(key == 11'b11110110000) ? 47'b00000101000100010010111010000101000111100000010 :
(key == 11'b11110110001) ? 47'b00000101000000001000101010000101000011010000110 :
(key == 11'b11110110010) ? 47'b00000100111011111110101010000100111111000001101 :
(key == 11'b11110110011) ? 47'b00000100110111110100110010000100111010110010101 :
(key == 11'b11110110100) ? 47'b00000100110011101011000010000100110110100011111 :
(key == 11'b11110110101) ? 47'b00000100101111100001011010000100110010010101010 :
(key == 11'b11110110110) ? 47'b00000100101011010111110010000100101110000110110 :
(key == 11'b11110110111) ? 47'b00000100100111001110011010000100101001111000101 :
(key == 11'b11110111000) ? 47'b00000100100011000101010010000100100101101010110 :
(key == 11'b11110111001) ? 47'b00000100011110111100001010000100100001011100111 :
(key == 11'b11110111010) ? 47'b00000100011010110011001010000100011101001111010 :
(key == 11'b11110111011) ? 47'b00000100010110101010010010000100011001000001111 :
(key == 11'b11110111100) ? 47'b00000100010010100001100010000100010100110100101 :
(key == 11'b11110111101) ? 47'b00000100001110011001000010000100010000100111110 :
(key == 11'b11110111110) ? 47'b00000100001010010000100010000100001100011010111 :
(key == 11'b11110111111) ? 47'b00000100000110001000001010000100001000001110010 :
(key == 11'b11111000000) ? 47'b00000100000010000000000010000100000100000010000 :
(key == 11'b11111000001) ? 47'b00000011111101110111111010000011111111110101110 :
(key == 11'b11111000010) ? 47'b00000011111001110000000010000011111011101001110 :
(key == 11'b11111000011) ? 47'b00000011110101101000010010000011110111011110000 :
(key == 11'b11111000100) ? 47'b00000011110001100000100010000011110011010010011 :
(key == 11'b11111000101) ? 47'b00000011101101011001000010000011101111000111000 :
(key == 11'b11111000110) ? 47'b00000011101001010001101010000011101010111011111 :
(key == 11'b11111000111) ? 47'b00000011100101001010010010000011100110110000110 :
(key == 11'b11111001000) ? 47'b00000011100001000011001010000011100010100110000 :
(key == 11'b11111001001) ? 47'b00000011011100111100001010000011011110011011011 :
(key == 11'b11111001010) ? 47'b00000011011000110101010010000011011010010001000 :
(key == 11'b11111001011) ? 47'b00000011010100101110100010000011010110000110111 :
(key == 11'b11111001100) ? 47'b00000011010000100111111010000011010001111100111 :
(key == 11'b11111001101) ? 47'b00000011001100100001011010000011001101110011000 :
(key == 11'b11111001110) ? 47'b00000011001000011011000010000011001001101001011 :
(key == 11'b11111001111) ? 47'b00000011000100010100110010000011000101100000000 :
(key == 11'b11111010000) ? 47'b00000011000000001110101010000011000001010110110 :
(key == 11'b11111010001) ? 47'b00000010111100001000110010000010111101001101111 :
(key == 11'b11111010010) ? 47'b00000010111000000010111010000010111001000101000 :
(key == 11'b11111010011) ? 47'b00000010110011111101001010000010110100111100011 :
(key == 11'b11111010100) ? 47'b00000010101111110111100010000010110000110011111 :
(key == 11'b11111010101) ? 47'b00000010101011110010001010000010101100101011110 :
(key == 11'b11111010110) ? 47'b00000010100111101100110010000010101000100011101 :
(key == 11'b11111010111) ? 47'b00000010100011100111100010000010100100011011110 :
(key == 11'b11111011000) ? 47'b00000010011111100010100010000010100000010100001 :
(key == 11'b11111011001) ? 47'b00000010011011011101100010000010011100001100101 :
(key == 11'b11111011010) ? 47'b00000010010111011000110010000010011000000101100 :
(key == 11'b11111011011) ? 47'b00000010010011010100000010000010010011111110011 :
(key == 11'b11111011100) ? 47'b00000010001111001111100010000010001111110111100 :
(key == 11'b11111011101) ? 47'b00000010001011001011000010000010001011110000110 :
(key == 11'b11111011110) ? 47'b00000010000111000110110010000010000111101010011 :
(key == 11'b11111011111) ? 47'b00000010000011000010100010000010000011100100000 :
(key == 11'b11111100000) ? 47'b00000001111110111110100010000001111111011110000 :
(key == 11'b11111100001) ? 47'b00000001111010111010101010000001111011011000001 :
(key == 11'b11111100010) ? 47'b00000001110110110110110010000001110111010010010 :
(key == 11'b11111100011) ? 47'b00000001110010110011001010000001110011001100111 :
(key == 11'b11111100100) ? 47'b00000001101110101111101010000001101111000111100 :
(key == 11'b11111100101) ? 47'b00000001101010101100001010000001101011000010011 :
(key == 11'b11111100110) ? 47'b00000001100110101000111010000001100110111101011 :
(key == 11'b11111100111) ? 47'b00000001100010100101110010000001100010111000110 :
(key == 11'b11111101000) ? 47'b00000001011110100010110010000001011110110100001 :
(key == 11'b11111101001) ? 47'b00000001011010011111111010000001011010101111111 :
(key == 11'b11111101010) ? 47'b00000001010110011101000010000001010110101011101 :
(key == 11'b11111101011) ? 47'b00000001010010011010011010000001010010100111101 :
(key == 11'b11111101100) ? 47'b00000001001110010111111010000001001110100011111 :
(key == 11'b11111101101) ? 47'b00000001001010010101100010000001001010100000010 :
(key == 11'b11111101110) ? 47'b00000001000110010011010010000001000110011100111 :
(key == 11'b11111101111) ? 47'b00000001000010010001001010000001000010011001101 :
(key == 11'b11111110000) ? 47'b00000000111110001111001010000000111110010110101 :
(key == 11'b11111110001) ? 47'b00000000111010001101001010000000111010010011110 :
(key == 11'b11111110010) ? 47'b00000000110110001011011010000000110110010001001 :
(key == 11'b11111110011) ? 47'b00000000110010001001110010000000110010001110101 :
(key == 11'b11111110100) ? 47'b00000000101110001000010010000000101110001100011 :
(key == 11'b11111110101) ? 47'b00000000101010000110111010000000101010001010010 :
(key == 11'b11111110110) ? 47'b00000000100110000101101010000000100110001000011 :
(key == 11'b11111110111) ? 47'b00000000100010000100100010000000100010000110110 :
(key == 11'b11111111000) ? 47'b00000000011110000011100010000000011110000101010 :
(key == 11'b11111111001) ? 47'b00000000011010000010101010000000011010000011111 :
(key == 11'b11111111010) ? 47'b00000000010110000001111010000000010110000010110 :
(key == 11'b11111111011) ? 47'b00000000010010000001010010000000010010000001111 :
(key == 11'b11111111100) ? 47'b00000000001110000000110010000000001110000001001 :
(key == 11'b11111111101) ? 47'b00000000001010000000011010000000001010000000100 :
(key == 11'b11111111110) ? 47'b00000000000110000000001010000000000110000000001 :
(key == 11'b11111111111) ? 47'b00000000000010000000000010000000000010000000000 : 47'd0;

endmodule

`default_nettype wire
